BZh91AY&SY�l>O �߀Ryc����߰����`�R�Z����   b��P((�$��4556��!�M4��A�hM�T� �I@hhd441 � �M21M0�&�F	���#C@%O�4<�d��0� dd�4�#��i�`��244$� 	�CH5OM�z��I�1���z���@dw( �~�h�D2$($u�n ��h}����� I~����ꊑ*9�$�M �
��H��9@�q�	$�qr���2H������+�f��׳^��i!$lj=�:nh���~t��n�ֻ
������.�pc��N���52:[�)tGI��/�$���[$�K���T��z��ѡ�+_Kj)�%;Nʥ�a����x�u��Z�s�1$#fu#��	St��0�=�^�i�ԅA�a�Vf�b��mEB�ӑԬ�gj%e-<Ơ�Y����G�a�\�z�6���"S;"��}!�Ŷȇ31��X���ݺ?*_	��OI�9"8@V��F(��P-P�a>��f5�'��clD\�\�1��I����fi�a���2k1����	����1���5��V����d�,z�˻�l��w�I +�>����[�ā-��V�H�1$�ؤkY�t�e7D7[z;C̠�� �BO��<���s��t�f����y��$$^Pm�#�
���*�E��a�5d�XI��V2�A�dxJ�����5�,Vz4���o�����	�}J}H{���/G����
�\`�L���?��t>�0`iE;������܏e�j���*Hʔ��^YD$��e&N�x���Lk�[7\:�����Ha}�|GL���m�h3�)��5�|}ݜѶ�������رh��.�@Z���)�-�(3�/(��[��!�NI�<��5��m̮�I�1��Z�=@o(*�f�5�4f^�؂bd�������h¸(;Zi�+E�%����1�Z��r��G�C�>7�Aȴբd�@��b6�E`j�Ƥ���!�q;��Y����f8-|��m|�����B�FK�q1 �d��!��F�_آy�l��∛�r\�e����U�n��Ȧ�<��J����Y�W^�ږ�d;��)�z���P�^��҇+��3kG�����m��1X��n.�6�-�0�M����������=�[r�����W�i~2�����K.5�W	�S�Z��|V��%�C�xg���z"��Yz+B��V��bM�1g*���7x:Ҝ�}�=
6��³�m�[��d�.�q�/Cƫv���d`�]�Z��uS X)�5�KM�$���5U�^��~��~���qdū�n�Q�=�e]�yαl�p��zء���7$8Ŷ�=��C��i�)L�3��y�������/g��Q����=f%���J/��C
.��U>�Z�/F7��ޖ1����+9��jnL�g.Ů3e��Ӱz�|eϒw���e�["��Ӌ(N���>q&�g^kqkٶĠ\&���Ve���rK�O��ڱ��4ĕ�N,^�:��]D�v����F��İѲc"�a����N��|����q%�4�e�Y Ȍx��ζ��2o��n��^w��\7�奙h[rwh�
�����~�5}H[��h�ϓ+}i�"�y?ѷS���N/ۂ�4�wG�>?�D�D�O��7�Y���؄����b��K�/u;��b[�R�m�^o*� h�i�4r����h�	)�҉�ܛԢ|��>+��B���6�5������b��Ib-��*v�NK&��Z��O�;��ͻ������5���"���M�+�m1TJ�ot!
�����:�3��>�$8U$�$�I"x�JQT�(�sTT����.��8�y%��J�*�ز]2�2ֳj[�$�JҽK/�X��VI%�)���Z��B��$!0�#��*�	�S�9�p����,�,�Ҕ�)3��?���ޔ*�(# ��+�tnpxg��~{e�',.���L����}�O�|���Ͼ�0���d�:����0_�f��R� ���t3@�N��o��D�|�E3zI� I#�,��t��ޑ# \� �8iUT��BB��{Ԟ�w/��pt����e�+?aՌ�'�����9s>C�N�կ̒G&�iK�A���s,��V�2�Y.����a���d�%�pZ��s�`pt]�*T�'
눈��T�K��6����t]IpZz��1�zt��*�����C�*f��z��!�!tR"��"��+k:k(F�m�`i̟��h��QSIJ��4�#�
�!,���O�!e�(vF�\��x���}���g;7e�����O�ATT�b���Y7�=u��8;/4���d��u�Q�'�]�<C���,���}��.��&������u�}�=*���CX�b�%��O_ș^嗯/0���LXxQ�ڛ�a`P�ب��s=��x��6)-�ai�RJ�DTN,XHJ�@��T���7��,�b�����b{.��.�`RD�qrZ�*��|B�'f��o��6��E�uÂ_PLbF4���(��%������=�����⨩���0_tA��4�*�F��A���6�_� =Y��N%�9���;�S���$��&���p�.=�	�'F�3�����QR�Q�۱@<�p}a�QR����R�����������b��N
`�@V�a{x��`��B�)&���Έc�1�y\>:5�I��z�i�ͥ�0���2,�.C/M�����3��՝QR��X���mq���(:��&уH�	|)��	��^4��A���Y��w�����dj� �|>Hv�(k�k�1H�5�X������#8b�:�#q�0K�Q�eN��R�j��V}�6$�8�=c$1���ܑN$%[��