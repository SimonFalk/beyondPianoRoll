BZh91AY&SYg,] 	�߀Py����߰����`	^{�i�  �猦�]�]5��	�PMꞢz~��4=A� z� 5O���hC@ h   �&L��L �0L�0�D��z��h4 �b 4�d  E&��<)�d���Q���=@�L#@4=L�D�	<��z�����i臠�� ����¨s�,�"�QȿS���8 �H~��CT!*�@R�-���bh*�(4�bTb���b��ȢI$k�Hs�Z�"?�H+v�qo��e��J ��k����팶�E��¢NG%Á��P�bb���V:�S�r�#Z+uN\T�rA��1Z�u��3�S=f�:^cq�6u��T�VR/'x��*r�la�+�QJDA����6�"��Ӡ��Ii���N/��$�4�I	�&R� �A�1��Mk�ssP*�I&�{K��~�\��9Q[�Z�{l�8mf�b$``��P�)���G�3T��TǃG5MʨN�
�t?2+�\>;�vS�B�O}���M�1 z ��6l���!�P�E��^���1h27��U0�QYDP3>""����00z��*O�4�r2�(�Y`��`-"�-м�'b�Lu�x�z�]LC5:�,q�^�|PJo��aPV�D^�~�Dx����^��@YB�yx��S��1�������;��5�����EF+n��ZP���bfY�_v��*7Ӏ����
ʅ��NYj�Iq�0T�+"n����Ͽ��:f zi�V�;èO�&�F=h���~p�WA�Ċ��cȓET��H��v7o�=t6W�[x��r�'|o�BE+�g��(���9~���A��85ͨ'��
z��h�h ��ˡ�8����r`�t��A�N&�9@��:�?2g�y�R뗮"���H���w"��8Y�32Ӑ�	X!h��]оtH��2pN�)VA�U���4���~� ���F<;dt��$P��-_Y2Ԍ��Qx��s���e���w�F��Tr�	<h9K�љ��n�����19��nē5�5I�\/Ȼ{��1}B��/,ٴ�s��v�2Ksd��qE�\�.Chi'��Q:��>�� |C�| �'h�m��� ���I$��cɅް�T��&��A�Q"L�$��lE���-sj"�BRp�6^�ɐ&	�Sb���La6���L���XP��LJ��> ��!�la���n~��0�)=5屣�_(tK�����Ȭ�<t�7��c�2����uG'������8bi�44��
�3א�z_�������"���y��X��H��l��|�A�|R���UM��	o�"V*Z:��B���y��c��݃�Ag�;���@G]�u����^Ty��d�
Bo������2�CH|D*��XA`�G��Bt�*5��\	\^�ŀMsI$�AV(�(��T��Ǥ(b�d��f�a6�*�"(	�X�?�Γ��5K$80 )E����.t��pSO��N���	�����T/��5�`�(�b�.w��RI$K�:��h'�ԗ�j�#<9uff�6H�=�U8��� b�i����jFôQ�Y��2dK�2�Cx��e���3�Z��mm���j�ZȵT(PW�5$� e����aJ�1���rl����H@�u���ހ|x���*����y.4�tٟ5X�8�,��b7���$�i��gd��r.L�-F�!A��Ϭq��"��� �=��UM�xyx�᰸�^ l��c�PQ"I���L�'MU��뺀����όPJ���0+�YIT	���l7�$�.=Z��δ�l�m2A�JY�ܧQ\{z��l0Kf��EJ��JP�� ��v�/e�����.[�[A��}J����K2���u�!РI��p�E���)��9b�