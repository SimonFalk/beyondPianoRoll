BZh91AY&SY9:d�Y߀ryc����߰����a,� XR���)@ (� @ $H�L�AJP��}���    �� �   � E�����U�P(�� ���)H�U @W>� �  x� 0v��ׯ'xe��^���t��7�v��=�+�ďL��!AP��}h��*�޷�4>��Tz�=4to��{�z����=i���z=���ޥ Sx T� �.�¯5ؘ5����Þ��^��k�I[�v�����۽�ݺ�܂��
Tܶn����yn��n���{�9.�&�u\�eݻ%ۺ����x��' = � 	��mV�����uX�m�ݷq�⻳�-/ON,��on��xJUQU�mA�����v�:��smcf��c]k�g���l�E<Q%J�   v�pvkӻu�ݚ�y���\z��{xKT{e9ۺ�n�&�w��`�z�H*QJ
�{^��{�쭽z<��vzz{��ii��1���vtyEQSp @�Jper�dק�-6�n����S��^��'v5�/{ӳz<v�RR�PP�=��7�/Wd�v��M���i�ٶu��k�ٮ��d>t@                         ���d�J�Dd14z��  �)��R�!�!�M�F�44Ѡ���5T�z�         jy�j�$�Q�h 0#F����h!	�T3Bd�d���#�ɂ�� B	��i���'���h�L��Onϑ�����|��?��g���n�h�3m���lΛla�{�m�nv��fm�f�?����7��������a�J��u�m�3m�pso>���p�]�oBOj�� ��x�����x��?G������v�������{��m���ڶ�(�����j�6հ(Ʀٌu�ãv���t���/w�y��^/o�����7��z���s��m���?7��������P�Wa!�N
f�9�v+ ��lSN�v�Sf%(���1�&@��6�e�Ls	X+��Wh֮��k�WI@e�ǆ
w���p,��ck7�Hni6�fb �R��p�6�.|�O
P���1�.F�j��ڛ �讅�+�L���s��F������7te�7f��/x[ϵ�q�}2�6q4�F$�Z�5n�a�r�[N�iq3�zA(*�˥���v���5�eN�Ϋ/����s);�1��6�Vj�9� �Gsb����b'��
�f�W�x�i��N��+��(%j���*����% ��.P��;�Yvv"�1y�q�L��z�eذ~�I�1+�``ɜ���7hn��}�9�&�k$1��,��`G���$Y�ln2-o�{�2�r-���>2�t�q�����QT��є0�X��(K'3�Z�sM�s��n��:��^]Њ�טi;�f�(�M��I#F-��n�V���j�y�Q�X���l-�cgq�[R��y�y�Z�eK���r�ͳ��A�
���������V����Њ�(��u�X�ѓ5��� ������̥V�;vc���7,��˼� 9nHl=�d�T�b�7QI�d����[��h�S�J��������&%`�)���,�&�uo-�
����O%��s&Sq9P)ʫ�1�6RT%�a���*�P�u{9��Պ�^���0;x+v�&ѭ�On���&]�q&%�/)����.�f�ZI��պ=�rG��}�O/����mis:-��yvz�����Q�]��˱�=���6����s(��s1���U�^K`��VXsP�S7!"fZR�Pj�I�Z3K�ok4�3,0���-���%�6�'���%� l��c�f`���d����չXw,�����.�m�s���`k[�^�T��޹A���Ӌ�����IV#��V�{uo_J���u|a���2�I�O!W�`�uՉ�֮��m���e�y�n��q]'�m r`��ޕ1^ݍ���1�&��`Ȥ&���C2]m�d[ȕ/kX
(wH��M���]�S(c9�[6�]	rc:,��q�5cmT2V�hV�s5n�7����x�"����	�b�T�ڤp�u�R��	��-5��M��p-�7nO�L��z�^�0�5�sI�[������R�	<.𣺙;i�p�ڡxDjF"�G�cs��ޑW�,��H#Mm껽��\l�0�n�e��^m@�x�l�hf٩�OK���J㗚d��S	ތ̔�������h0���w�N�	�2��Z{\���~����7���R]^�ѦM����Gp���l�ǆ�b��5�]L�*�5BB�����>�����%]J�\���	3{������x��@�e��6��ʑ��z�ͳ7d�H�]ܛ.f�5n=�M\4�L 7��tm�Ƌw��N$�6m��0T5��H���ǚ&��b9.A��`<uyӓ���s&g�ނoDTL�D �@ң��]˗����ks��Y�%IF�*rS�g,��'$g "Qדu�t��Yx7.e+"�r��l���+*Z�5-�/"�8
T�[W�d�6�v�VH�".*ݰu��5!�t�f���rʽ�j�&lڅ��8���YcA�jM�;B�p�j��՜�V��tT����}p�]�
��ofeH�[��-ٔP�X�p�
V\���;F,7����H�Dͭ�V�-�4'4�5.�6e�(;7k-�L�%*�k4��~:I�e���@�HN"�,��t*�0�cm$ꐄ�F-+l�/(��,!�_Z��TW\J�����E�6ܰ���eҽ�,��
5�0/]�lLѓq$t�qPb�RօI�2�G{Ǳ���2�"��U1�f��<"b������*�[y{�7�VQ(�6T/2��y�t��'v�3J,k[d2�(NL��'�[��[GK5D���6�$�Kp@�e��!��̚I+�`�5��T�H���8a�zq�z��<�nL�B��#4�kooh�޷L|�4���b,(�Fb�@�3b����SE'�^h/*MԹ�P1L%	��H�Q ��8q��Uwq%�����ʀ����ݵ�lڈ�ot\ܔ��mKɑ-���@�TtJ`T\�I�{�1�&<ô�PVb��Ut�u��F%]&�7V�'�M�aĉT�*���v\d�b�b����mS���&�/���RV��mmɲ��P�5J��3*̣N�n�n�nؚ2�dʉ*:F憲�nc�_�4�a�**,��
�Fa���N�՘ �`Ȗ!K<rq�����Y�^��R��'V��U�c���v�Z���L�o(H�1��
�y7]����I㵘�к�Qm̱�k:܁�r�cqg����F�ƙv�K��M�M�ɧ6�$镊JU��9fqY���dr�a����K���kuؽKC�;lA����bj�	��dܡX���E�"���aPO7�P標c�Ruַ�ݘi>�W��V��t�#����׭dkl�,k��Q�����6��Z/74̜dUiފ,k9Ic���,�F�x�%�s��B�F�DoYV��:�rѽ�+vK9�)]���><9� �܎��Ae}-fK�N1�j�Vs1�%5IU�:5�l�����g�rn�h�T��t�N*Wj�X�g6C!Tz�sR��u����&S��C�1�dtCNuY�A�`�9�eU��P��V�,��V#���h�)���W�0e3m�W
w\��@���q$x�íU��I\�ZP�\�x��+�T����{���\��
�][0k�"�=���:���G�j�dM:���^^p��L�8i�ǵ�2���JZ ����,^��a�3N��OX�m�xS�j�%1AZb�F�_NS�tu���c/Lk,��p[z�qX�i��^@S��;�ݭ�e����C.�)�ɬ�"�p>]o[�(=�l�����n�H�͕tͬ�7(��f(�H��3)�
1N&�)Q)�*�LK���3[�Cm���&gd4��YW�9�+~S�$�Tb��U�k�r�rxt�CzehTNܱ�_�x]���E�qL�F���gb�gm�!s����P�����.�Z�!�%<�zѡsd��(���5�c��n�8p����U륫*�4�w�Q���RZ����c"��z�AXRV4̀]l�\Ë]+�1�ctY:aWR�ʋ`Tݐ�[m��.O+�kO$\c*/E9�.��z����Rb	���]�`�G*k�UF�f���ظSr�W�M3z��y�?�7D\k�0��@�F�h��3	&a�Z����4.��	w��>Y�$ʛM��0-���mGO���9���<��P���xA/�o0��S\��Y�q���JD�G!dm�n�����{6��ɋ-�D)ws[@����8��������/����O����5��c����w�ï���׻^\g#��t|W��S���$�?�3Jq|.<f���+\t�Ct�*�b{+a�:����M�0�8֮k�bn�5�ڸ4��b�ˮnDѣ����<]R���O\��8��=��k�y�5m����q�e�G(v�w:�a{��pk�n��1��[�3"�D�c���`��8�tv�tq�(�e��uͰ<[�ۭڣIm3�������u']�0]�v�s�Շ��Y��c���x���;��y���Ѯ���xy0n�.akpS�E�%����d�o�=3q��n,�n�����]� �tq�vػX����;[\�Z�a�M�W���
<,�<�lv�8��.����6�ձ�fh%�;�2\Y�/��̖��k�m=�6�;2ݎ��z�{�u�T$)G��r<�Cw�)��CA�'[%�uv�:�n���ݞ�p�F���E��!�Ʈ&�m�w��Z�,s�_�z;���uù����֮&/�4v8�ch�D��^ݔ�Ś�;�,&��E�)�n�l�/kf�oX.�����H�����[���4�ve띱�|c�Y=�rIYK�ۜ���M�q�r��Gk����M���=vwF�+9�α`��r�&`ݷYw^ݹ물�k���<��O��<��>3��n7&�6�펶�&�D�DCn�8��G`�ź{�9�6��7���3P�e3�Vm�N��wv�\�c�����!��#����=1�vq�=o��f-e�/j5'[U䄯0�0QX��Z�݈d6�AI炵����mZ��nZ�غ��f�܏aNz$�mն�WD���v��77\��:��[��R8m��s�ոu��3��fB�����n|��+Χ�[v�^v��zi㎏;�N2u�]��tx���1�>�ք����pQG  5R��T��-�����5��f��ͣ����{:nxm�m$��6r��kv�vʣ�s����Z�:g�XB�p�ʸ0�P|=��؊W�25Ɯ&��</h,-��Z��V�!�1�'�)�rb6�%�c�!j�
Jb���cL����lv�[3eRCX�H� V�rM�v��ώ�:,��s��9Jn�p+�XoY��u���o]'L�0�ф���g1�����,u�ۂ_͚�δlE]�'Q�mϚ���'0M����7s�Y� ˶M׳۱j�kq��u�Oh���vØ#��ݻ#ڵ��r$G]��9f�W��Rm��9ƴ˛��i��u�'Zʢ�Шc�v�wh�A�s���j9��9���p��a��X�Gm�bdv^�V�@n�.�j�ݮ�Dc�mn��s�ی��+�bmvSs���Ѥ���嵎;k�v��=��G�Y�����\TD`���GSD�,V!��O�d�n�㭼��j�0���*r=�M��c�6�</�Q"g�v�`� ��z�wv<��6#�����h,�������瑜���ŷ]^�=nu'�ᣯ=��a�#�Gc<tb�u���sd�=��ĺ5�m��c��]���[�ڞ�uj���6��7$e��g]��y����OO��E��خ�]��^��U��ۉ�{�#3k�����a~�{���,�s2�p�b�v��PЅ�k8���4��]us�j�i�d��_r?3��n�F"ݍ���v��2;u��}�����9n���n�X�u��N���������Rytf�Ǐ%Dۺ�7&���3��ӝ/$�	˨��_���Gj��:�ɣsX���[�pc��M�e�5�6M����c�L���Z؋�Z���.������:��I���wC��f��kdD7ls�2��wk����_=��,Ck]>��\�����j��is�����b�,3�-�vv��8��n��G�GG!����YKt?Vf2�jm�z�Њ�NrY=\C۲�m�u����+X�Vp�����V����
<)ƵӉZ�X�8�]�ɓj��ܧc����X�V-�U���m�a�lum�XKl �ֺ�=u�"ɕ��s��������l�1mj���nm���i��8D��W\:f&���ض��w�i.��s�=�2z-�ۘ�{s؋l���B=��S���=b�.W���Q���z��mӁm����o[9�[t��=��(j����Pӝ����6t�F<�6��v�sf�{]�l�@��g��\�Ø��`�qu\n�s�x�e1
�GWֳ�+��F�,��6��7r89Zj��\�C�G�׎�.��ʕ]��[6�bx���$��u�l�NM9@�$C��:�7F\��㎊gƸ�Cc]5֫r�!���Ԯ7A�!�v�*:����m�Ȯ�n��"+A��l�at�^sp<tTseά����Q�*��]v�`�Xz�E�u�S����Wۣu6�]�o9l,!����A���u[uM*ƫ���k���X����Б�α�Ε�-�\�e�Cb#��vt����8�Wgv�����`8���Uv��b�rp�p�����w3�M5y���ؾ.w�}�m����u��y{;͛n�u���;����6�Ǐ���{_��UK�~�����`??_����ެ%�4�k[u6Z��X2*�pA�n�L��,5��W:�m�+��`�Հ�uj�R��9k��ݤ��T�o{���`�s�B�0�;Fh���9�$�L�z�uNn��Xl(�����q���!���Q�$Ѳ��ToZ�;^�	���0��!U#��*t3��̻�<���N�m�621|�d�{���6ݟQ�:�*rJ�-�_��Һ=�B�����W��д���J3�fR,/Y�ԼSYs�f�V�F���w{Kg�q�J�v��l{��<��A�&�w2wc�5r�s<�K��5 ؑ������[�(��5���u��cs򕺃Ԕ�Yk�����C�9M]α�N�-)�^P*���Ô�Q=�Z�3��fq��8�<f����Ui;Y۹1j��FMU���]�5bM��te;2��3(��;�ϒ�k޽yV-�e]��"=�ɮh�[�B�ʧ��#�S��.�E�Bl��OK[�ƫr��z`(�,����W�]:�j��VV�cU����0����n�b�aP��[E�M.�c�a=��mĻ��Y��5,f�*�t��}W��8�\���yFooZ�z��d�s�Q����k4ֽ�%uZ���S�ޥM�1q�����\�1Ź�97���aa�#p]\����Ԇ��μ��2\�1B���lA�˧Tl(�M9Z0<��Q�wv�wK7VfpC4��9l"�Wr���]K��Q��e�oK4c2�pk\3u�2_4u��'��e��{0�o�ݷC��o�cB�݆�u��6��3!	bb��KG�-&{�?xr��i�)Z#��5�V�o#V4���1��u�Eiʽԕ	;�a��}���2�(6v:Т�V�L�ɏj4�S5�0�,�fqV-��/"����j�����k�R�[�f�ś9�*�h��0'��� ���9#O���Uv(f.�q��w�s7x�j<U��k�6�f�`v��P��;�{.t.�o	{2�[[.
k�����O5'-�3����	/�f�t,��?K�Ӝ^!�c� ����}(S�H\�j��674 f�ۅrl����n��N�<y��9kk2��JdNkA��j��y���*.��РͶ�a���Ӯ�L�yG/V=��n�aU}���r�[;��؁��z�6���R��)!���e�RĮ�x0]o_U�e����4S�2��z6��KE��K����E��;��Hc�,��Z�g3gSD�&a�����F���څ���'��$A
�Q�D*Mh�M;�n�?\�p�:4��gm�\J���0,T�{��]#&�|{���V�F`�F���uӭ�o7-�ݹ�� C�̬7����.��x�y7{��b���稲��i��]�ҙ�'&4�zm��M�WM�ZD:��`}3�D����b���T͗Z�e��v}�F�w-]ΈD�Y:���p��ʲ.���.��붆uv=��� v>�/�c�{3�ݾDvl��a�=�����<�bM�:�4�V��+m��FK�#k	��\8����w�	v(�H��{����ʽ��np[����1ve�]���^�r�`���1@�33S{��z�����W��������-ʕ���ZJ��?��˘9�[f����=d������(<�NcQr��@�N|�9q�k�v����L���N�x��c*���ӡ9Ɯ��M����,��Zx(�t��5�^5�A[����s��cL�l<U}7��Zln�G34�H���1�ە�֪[V�7�^ay㤆N���� +-_ǻu:��痥�P�6�ڰn�D���]B��*<��)�)��ИbE���uӧ��h�y¶��b`�҂՗�s3D��X&p���anR;]��.mY�'F�� ��go��3rv��/�����(ݛ��uX7��U국�#Bj�����јo�����wq̻6
�pwH�[�F>�Won��˶�;� ��v9�,z�*ӌl�T+qaQ��maNMWgq�A��K+�PX�0'�w�H�PX 6o4@Z��sFi���4"V�-�R�-�Mv��-u�&=������y����j}�[�o�h���%�3��YۇS۔�[�(0�+q��=}���e�@�̚Q��v[���(.��jxNY�\�W����U�M�A�2q�P�ȓֲ�ܙyo�ER��C���7׫���V7Uf,!¯�j�8�ed�p���qa���@��gdķ�l�՜s�X�j����v�;��E�/��^u�9��"mu�,'Ԟ���M����H�+'n'&4��:m��nn`���f�{v��ږ0XH�v�c/K�RSf�b�!�*`���R�M��u���h���Wf�t�v�h"cV<��f ��`��[R"����k]+�]�*Rn�Q���,��뗚3)�A�ZR�!�����\�TdkȥN�;{71U�3^�چ$�2���yoh�S�m�!^�J�ԩ�T�-;���oXY�
��V|U%iP�nt�-�z��5���am�����shƵY��5Nh�*+�m��s���s%���3-��V!8�f����>��L�R%� ���[NGܺ`�H|���]n�����}{[�*�xᴤ�\�Y�[����ʈ�p�x�-�F��E�0K��FeK�k�ma�,񎰋��]��4v�g�.���@��bLݜ��sP�.��+oz͸&g(%]��+,�f��ˍ�Gdv �����(��q�3v>�t�Ԩ�|�=k&������0�Fm�	��Ď|�>�.aW�H��*�����Y���۹4P6��\�햶s/CRU�T	��"���[8�Y��.�"�)�D�L�
��Q�u��Q��$�D���#�u�d��	�du�˾5���v�T��ZLb���2p�oJ�4��x3y�<ŝ]�ZV�����in&o�M��e)De=��GỦc�S�0��,`�'1S�9����Ծ{q��o���ɧ��m�Z��Ni���*���_i�ӂ:����{m�R���� ���kk=o'7\ӱ��`����z�&7:��zPH�?^4����b8.$�uԓ�&ݗv�\�K��r��5AbL��v��)u$+��Z�U��Cc�6`�ѩ:�񧓧v����g�yA3abVηC��O4��61���5g,bTU6���@nԧ�����X�Vj,6Ɠ5՜#�|z-�U�>��o�^�\7TX֨�+�A7&܀�{2�B�+��i���T!����x�`ƫ�vO�0G�ۃd�M|9{x�p"ן�<OvU��m){��NvN�Nۆ�|7�;#��a6,hK5nt�
��5��1X�݌n���mE�������-�pF�NC��_C3���t���<8�W]��L��36։	_���~N8���q��w���wM��O�@���v�B b�,�]������ػp���ŗ��:Ś��ϫ����B%�v�z��	(�l�4��N��ӇE);l�[F��Q������7Mu�uV�[zŷK�A�\\�Gm��I�!q<��m�	��<å���1�����p�Mؗ��=�yc��6퍃vK��n����4#�:|=q��#u�����oZn6'��N�ą��SP@4�0��paUCB�mP�
6P�`�u�ݻrH��z�$]���^^�s	{u�.{Vݹ:Ƀn*履��'�:��n{'��%]��s�Y��-nI6���v#���w/l-θ�]m�$�og5�k���آe]�i��y���]��:^�6:�d��]�.'m�l�G�"왙�]ś��l��k�kqs��n,�<ڲ\֫���n}�=q��ݹWF����H4k��v��mG��,����������q�4	F�ɬdݷVѝ���jKOc�+���dڎ��'�X�d�8&�[�&y7&�(�8�_;�곌Zٟ�۷A鳴f�wϜ�&M�(fk�	V���]H���L{��Z.�^kڐ��{���ؚ�4ç-{�76�;��;�آ1���4�L���]m�L�y�Nؠ{P�%��V]�y����?yF��D��%��$�\�d�Mnb�3��:���oS\��Ɏ�'.�i���%i�uʞx�}�\�2=���رW��W}�ע��������93����%��5�DF!�HV��v: en���c��xk>��)҄v�r�b�f��c}FmI7�E4�+ ��;���jP=�Sj��3������t��9֘��Y-9L=�ɛG��ﾡud��m{�W�����Y`x4���B4����Cb��+t�;]]�]����y{k�E�%u�h�WG'r�&��ev�݀��c<F�W�A0("J:�r�R4۝Rfhagzg��X���0]����tvX��>t@���q�M7a��	��'q+%~���ӓ�hG���_7|�kT��~��S��c�)�.`+�q�  �UƔ�N{#�x!|�f�g �Q�2�$�}�mùD����Y���!M�N� �S�6b���Ģ>m[��3#m�2������?9�Y���G�n�Ge$D�M�z-����f��ҪD�ҏ���HRoi-�l�����%Y8�j/�ѧ�f��T���Xz�+�.XQ��s`�*���ƣ+���PÖ.��C��P����	�X�B0��A�q���T	$��Jȑ�X���j��>��p@����{n?7]M���Z�&F2�&)��aK�麗�v˗�ĊIzA_b�r�n�ϼу��<��/��1 ]@���	�J��d�p��:���"9������` �K�S]!�i�pD�VK�D����\fvm�[�0�9Cd�qچL�b
���>��c�f9"����`��>d+���嘻}�i����R��ky��w	��I��b�l���o�{�09V��p�/Ri�#s)OG�R�#�pU�S���2��]t��&��Y?q��	0�"�����}�(�4� }&�$���}V���Ґ� 0U��Ԉ� e�(!Nά/��o���B��	g���=����3�L4�'TC*�V�t�+Tk��J13%��Ui�X�_V©��p��aH����S�7��E�q��l�M�a�B'��[�լ��h�G��:����?|���f�b�H�Y�� s��,�Ϭy?��c�"<��~�����:�Ȇ�@�?w�lI;#BL>�v�i����牶��t\�흳۳���������]aWƍ��p�E��,Oj֋�fL�s�f :+��G�ʖf!��V)J�銭��YFA&;W<����~SAÌx5QJ�%;RA���M���Sb-���s�"��i�TDە����␉�0���������ٸ��_�Lhm�jw#��P�7i_t 0?�s�*c�c)�u����şg$�	Хj�௛��=d��
�G�h%P;� �D-��'�=�4���I6���!8�6�>%�;*�;��p9�O�1�{��*4����H4��� :�P�C��M��*bѤ�k�xW�2��9��3���u%*G&X��" ���;p�s�j ���6!��;b�4�>��uF����@
��Մ��:;�$�x=�ԏd3�}�L8;�]r$�RF��=k�<�wN���^��4e��B�8�n@��ې���;��Uw�e����琭��
い[�{�~��"���>GѴ 岾�g��{LW�|�K�w'�R���K%; 0
D�"�H��J�
 
�ɋ�f��l�M}S�-5�2��r1�~����]���3�d�'ɴ�����1�(��������.��v~?>k;�6xˁ���ʋ&G[���l�Ȋ��5�Ƕ�Vi��*y"	���u�q�!��H��I�5*X�+�
@���.UO�`N� )�%�`��ժ�rr>���.4=�����r�Ă���ZnV�,bQh9Qy?����%���0������U�.�8�u�5��-jn�)c`Эp�i*r��I-u�nm�E������������0t@~��<uŏbM����AB,�������c7?/*����p�R�c�xW�Hc"��p%+��x������`v�<Ȯ2;�)|�c�u���y�
):eP����s�)�V�`�����(�5����M�bG��z�;.s���)�������y�lR�[�칬v�s[];�k\v0^G���P�ȴT� QШ���z�s�zωe���_'�t��:ټ���fT��ˌ�.��V��j@aU��� ���:\����+\��;�%���gY0�ڀ���qE�`���P��R$|'�<�g�P(��k���*c�QX~�Y��mB�� �9��f�����u 6��E�J⡪<P�1��xŹ�`�c��E�wS����A��\�(6v�~��#�~"�ñ�4~�����v�=�v�)���i������`��uH�}��ȋ@��+B�|�^�߲�B
=��?��9֌Xi��,@�Gܠ3SQ2FG���GD&Hp'���X�a��1��϶N�9\�-I�jc$D���X�C�-�g�)Ҟ�$ �6�Eb�jn뇡-#���d���F�*4g�7���~���d���g�ߖ��7'.��7y	�S	r��F]�Z�C��1Cyx��O��<�`d�YK,I9����
��B�\�W��+	��QٛnOe���:����+S�����c��!)���R��6DeRV������k��om���eH\]Ry�ɞ�}x�������vZ\�u�:�c�ۤ��������Z+~A����K%��ǫ��P]���G����z�1��>ž�$�D�����{�<��mi46�_oM�U}�|�ۢ5�q�7peT$�5}�E�H5b;w��8.�k8!Sfm!��%�,��Ta���t���չY}���3���w׌�*�6�وɽ|��a�B�y�O���E\��Ɲ���&��u ,ꇂ3*j��SꙞ�XDc*J�߄G�Z�_ B��Zws�D��.	����S{.7l]*�B�ۡIӽ�m&��n�JHl��IREh���ۑG1^�5T��2��� 6q%Vϳt��Egj�^�݂2�$����4�@�b2�fҩS|�j��&4]�����`�k4���x��r��>�R�sΕ�e)�o\ڜ�u��ޖ-�2a�oN�Wu:�m��������y��jˠ����z*Fn֍L�̛I��
�,=�N)}1<��em�M�0]��nM�bC�N�����ة������m8J:8&f5%f�2�bb�<��Mq�7B�fT��;+k���ov�o��k`�H�8����6��f�o����e�-�h�J�g	�`"�A#':��TLW��n޺�3�3&˼�ym
t�@  �H �&zBD�޲b qN8$� �$g�|���)�>�f�:C˿�V�_ONY�m�K �D"y�JC9�xUئC����8��-�>l$QG�d��  ��d }Sx���D�i5TRT[��Tv�^!��8��]�`T`�@߽"��T�!�yۃ��jJ[�g_>�������椔,��q �� �0�	"�Y 4@�d�@��F�$� ���H�8�I���A$D oEw���BJ����3��;��j�㊗���i�z���s�' �9��U:VHq�Fqq�RV����9����#��v��!H�	D�;�:�O���O�!��8X�߯;����� �$L���x&`����,c]�D�n[����U"R$�A��|�ĥa�� b ��� @��  �n� �S @���H>���*�l:*��P8àЧT(s��( �I+ī2���T��$� <�-=�A1oX�M ��� $O�d�D�D����A`.�\�V<zq��]\ҪT5��@���E Ϥ �a"�` Hf����AdTd���d��1��:�.9�%(۷�.q����ۘ����Dn�% :iu�Y ?�9�&��ǗN�P�u�'q,�o�}�w��Tu`��qyOv���X��H�-�-H��`�����h y�Q�0"q4I�U�����D �-�^{�P7UB�j��g��S�=�dZչxګ#�۞^v�>#��'����u�[�k��&�j�������;��I�Hx{=V:_I��M��tk;7-�4R�,���m�g?������:�Kl��iH�2e
�:�ޔ�Z����^�-�ݩ�@h�v�!ۮյ���߱���(�� �WPD�� ?���� �$��@	Hs7�O�)V��8�6�޳ψ�IJ$�F�,o��l�~�o�ˇU*mM���r���E]�L@ 7�b  @��r8��A�߁��yv�c�;@������M܇��E�R(��P R${��1) E�L��}B �i�>� D- R �o�'��)�	 G��"=�i$�	�@u�D�� E�I�d � �=O����[�t�v766�(�Ky�R
�( -4���b�F	�A+�	 F[ �@5�A�l"�@"IH}�H���'Z�]`���}톖Vx_���CQ"����7� v>�;�F�K#,�n6͚���ʩ�&^!��-j�Р�ܖ��w}c�*V}�>��
g������Yz9痋�R o�c: �g l @�m�I��'[jN�m����� 
@�⯊�,�n�'$)��������[7>��m�;p�m� m��	9�@H	Ώ�t���#��H���L�	 ;�@�@9�JG>d�#��j���(�烳�u7\��'�pZ���SM�`!UB
@��f �BIV�>�oN�WG��+�x������U�� �l�4V� �o8qgͱv��g0�}x9�~7�*���@�|��A�U�A)�0	��X�.��� b�@�:�(ju�}�Y�&��;�3�x��`��_w�U��Ɋ�(�,q�	"�H$ �Ϡ�$_d ���s�9�U��w�Z����&���ہ���ӗ4�,� u�@?=^�BFI�I��@�d;m�L��� R sY �8����H��o~�{�t�<n�6��M��=�~�8�U��UJV.��	>� s'ȃHz�Y�$) G���M�Aw7��n���U�	)�Ɂ BD�\�9�ޝx͝<r崔�̧�o�ж�I#1$����X�\��aW���a��<� $>X�"F�ϛ�R��
�Z���@$�|�D|� 
D��"tlR1�),0�#�W��*^�|�#������>\y�5f���ؽ���ï0�0�,A������ 7�I���ŏ��%`]�q ��\(ca |� DD�� 	���;{ϣi<-�Rp�v����V6
.�^<UY2�L�`�ׅ���鄰<%�D�@��>6ZH�R �BH^���%ئZ�1y�D�7�'��A)��2�( �i�WC�2� 5��H/�>ݣI �	�'R f�IH����I�S���@��J�g��.L��ۃ9��ӌ��88�@}P�@Do|��Jm���ۋoK��*#�9gu��nP z��@��L�s8,>E|ơ^�ʟw ������s��sԂ�5:ӲYs�-��m%F����R�q���=�m�ݴ�����AkWs��B=Mɸ��۳�ۂ�v�:7]�맵s��B�75gq����X��y[���bG������%T@�mۗ��M�sQ��kAQ�j��4rs[��JI3��N�Gb����A�R��`��n:_��$@�|��H��� )} B�h N�Z��13೶�Uf� @����g���l�Ͽ�:���us+ �H��{g��.�C���;� ��-��I�؁$��Nl�$A��'^'�RY�bD�;�H/"ٰD�dA$ �H@	yoZ�S�b�@�@l�� h���(A:�� 7�@HH}��" ���M4�(܉�ԅhG�t\lb�㾾w�w$UO2*YQ�i n�H�;P��ӎ���JR�)��9�n�"��}J�J�.��A� �z��|��H��s��A�&>����h|�id3�:��.`�6v q�S���IGU��ǈJ��9���w3�@�J@e0Du���&�I �$y�=I��u 6�D}��@�Nd�� �� �Y܂ BC۝�r�:�m�3�:m�1k R �{��@͐ /�DR!$*@�@R+��j��*T!"Gu��	#��܂F��b_X""<�����&�J�TA�!N�i�WU��W[I��l�ZU�ag!�"@�� 	�0LD��>`�$gΐ4�3�Z��F& �IH����I��	H��d��rHHH�(H ��C�x+�L8�8�{hx���W�D�P��Lon>@�M��㲤��蜬|e�w]����r��'��&끻v��S�!wSPHb�3�B HW"���V%�@f�T�g�Ҵ HϪI�`�r 8�����;QбV�" ��)|vDB��4��2b��a�\�Z�;�����v�v1ժ(�:�
t�A"�7e�6-����@
|���o,�H��A !!�Ի�N���$b'�3��I"� 4�;zs����<��w靔�Վ�u���j]ʄ4�Y�0@�Ag���I$�	l�dD@�od�R�UC��p��HAH�u b&�����z�<�;����s�r��>D��u��ƢO��wF�|M������jbTӎ�w���X�F��&�3��{�4 �v!Phu�"��!�0bn�4�?d���]���D7U��{<�{n`�R�-�;����}IRK�@�@��D��|�  ��
�<�H:b��3��sE/�F G��4�@�H	H�X"�"[�v�>o�誝K�g y� ��0D��J��� k�@) w�>�i@�܄y ���@j� �M��H��@�h�BK��j����PZkMo�?m�o��k���m�T�68��}W�[�b��s�[���8�=�e�
E���e�22��,���ajey�(����%���ɝ�U��'Y�hLt�8�rdź&'�Ӗ&!sN0�4��SBx�UC�&��=�D������5��g݇i_Ih|�2�""��;f��ҋw!SC_n�E�T;A�J�[{��n��1���Ί\��:�^K��j�^=�r����L�,+v�؊Htcw����qZ���	������d�7�ϭ+����M�y�̝����ɯz���<2�^�X��Ǔkt�@Il�=	��V�H5.�Gz$p�du{�b�?g��5�\�^���I�t*�NX�}��e�Gm����y�Br��%�+��+�љY�;�F{�.ɗwㄒ����{d'�z�bwKCη�\�+�{�\_n355EܭVA��Sy��=�Xy������~?=u����]���!�Z�Y��7��t�0�k�g9Cn{�j�]`5�$y�����F�mcou�M�|�=����n�*��8	�{y����i5� 9e��ewk\5v�/[�:���
���qѱlOa8�oGF�suέ��v��ݎ�[mgt�tV��r�;h��ԝ#�j�9�V��k*���0oj֮lQrRɷm���8�����e��E5ț�d�}���o��meR��Æչ�\��s�u��'1���=��z�vۙ�g=h�;u�\k�;e�۠:���7�/F��
(�<2GE@��s*�K��{M�cU���oYc�[�!�j"V���(#M����Σ���y�9xN)��K���k�A.��[x�#���{�g����ƶ���fqƃ��h��v��Uɤ,u6�/pۭۛ��a^-`����&�G5�i�0��.���y����n���\nx��R�N
�����u�?HjP�"���bm+�e��K��k�d�G(F�-��Wo3k�.��Sn�
�m(.̝wV����l���C����Qj�n�D7�B��m&b�i�)�<Y���Э�[)�n*�U��V.��W���Ӷ�71g>Τ�,���ȹ��y�VRDw�3#H�:Mm�ޛ�l��x������n��b���Žy�z����Vf���93W%z��^j�m�xi�Jp�sz���w��Gao�L]���ŷV;{]�כf����D�q�ݲ0n�]��F��?n���:���!��p�vkt���@0��.j��:J�1��c���
Af��.^l�@�me�Kۀ�*�5�횴*藒T��6��.6��YyuX��9���mıX�W�&[�]Y-�W+�r��g����=���W9熧�xc4�u�n84�:,N����$�N&�d$i��Ĝk<��s�gD�w�"��[�'F-tJ5n��X�V��έ9�o/N��n*��ƿ&��;GFe[E��p�q�o^x|��C)���W>����@l��h�1z��CHx�s��RS�I�	w��q�1"��ڔ�} 
�q}�2�'��9A6�^�z���
"��x쉧�CM\uo��L�_z�_���"��-}@D)�\��|�	�<���U�`�r�m�X�j��33t�D�D�s�E��V�zQ��Gā������ta�	����4I~�0B@s�B��H�H�De�-���z��4�%���UI�2�o�9Zؖ%ƣ�]{���T��8���4�����GJ<�=��Uy�q���_���v��*���|a-7�yH^2M�7��<��zц��}�I���#��O��ℶ�%I�id A�
'k��8�Sǚ[x�iWUud��3I}�޾�Y#@��sN*��sf|��PHw�Vm
�rJ��Ch�a'v�}�Dgg+� �F�!  �̻c��W��`�F�R;J^v�܊[%K���1�FO��}2<i2 8��� ��c�����$N�F�q��_��	w�
��ȇ��[�C	��������(�;2�8���Vm�Ћ8��5��O9".-��%a�D� Cx�=a�6Ti٧�A�u�ܼk��ks馐�}���Q�fSk�:�B� Hf�{��D$$�|�;�Gu��ԭN�<�XCf�:��YW�Q!&�6Z�>��F�O<�j#V/#�\���@
\����#�F��Y��F�����
��{�w[g0�����anˁ��oo�'�]�9|K��"��\��2$|DZB|���D=�1h���m��qB�RX�q
�җxm`�W*�f���X�H��� $�b%rj2�1G7D�!7�	�}��堋�����G�O޵��r�,���!O��2E��"��NIC)���1�v��ڪA�A">|Q{�kmD��V�� � 3�B�`�W���P�X?#">�U!	yH����V�n�R���j������&�Ϭ]�]��ʧ!�\rn������j��x��ۼ�j�Xӝ	�u����|�^;nT��+��s��EV�bT+X��$�Ume�8~w���W5���7>�ݛk���{�t�CF���X1�qp^� ������	m��즶B�� �X��N�	/?�B���H'l�R!"��Usz�*m؋{.�i^I���R���7�8Z�6O�#U�ϨkrD�-���O����>ڬ���@Y A�H̏^�M�j�� p�l����d\�3=�y ���CmI�*�Pb-@�b$f -4�|�*�RQ�H>�!�/U
�#�Z�"��Ԅ7w� ��ˈ��?S�"�\��
��ѥ� w��H��(�,i�+{M�N�N�R�f9������SX��yn��Ԉ�9�3x��Y�Ț����,ʇܱ��T�|�#3�`�ê�y��T	m��GQ޻ϔk�I��vE1��>fO�^C�Ů��C��z���n���մ[s��3��
v�
��ķ���T̓5�h�D����É����&�#袉�vi#�q��.7�N��5���I~#&�� ? ����H� >�����+ݙ�Uӓwpvf��X%8�YR����sE& �jB�[��fAR��Z��w�}�-e�}��sg�:Q�l��G����$OT#���W=�n_Y��N�#�nڂ�ǭLΔ�r�o�[��l�M��R�
6v!��{��[�.���1&��3�z� ~~�����pd�qV�,�����w�������Ԛ�xs��y�zi�0��_X	� Dz��6��`�q�� �4l��eS��42����*�x����� gγ8�C�gvs��]�� 9�(�.� ���ݻ��)�2��[ߦ����|��T뇅a,�9��d�Y\�z��8�Bj�$ᙫ�(�$v�=w��z]a�$�(�K�8H_d��<�N0Z�.=򁈦s��'s޻��w�%�8�ם9����\*�.�w+��sqO}}���D�U�Dp�"7!��ԕ��0���l��T���CȖ��S�'b�䊹Ux�V;ebb�K�������=sIQ=Z:K��-�B�7�8ݔ��pƴ����[�2�1�*$�j+0*JY��g*%k�v��S�ApgDKcvPC��ݓ�	R�F�!��T�HE�2m���yf�J�Τ��su��Y��ﻖ�n�wv�FG�����?Ac2�-������g�~y�8��cϏ视]�.�_#H��
�QFuS >�4,���78�Ȁ�A.7�t������Ǫ����<t�6��%�������:H�o䤟d?!!����of����	�����]�nޞ.+��m_]�!Ҥ��G���l��Kc�8@�{a�S~�N+秳�DN0Z W�W"�_Y}`�7QG����خ9�0�|Ç-
˴.iۺ��ƍ�1���c8�H֯�@��w�Cl�Uؑ3q���Q��W%2��Ya�t"!�R5t���h�0����z�xz��4�:y�]��'�ߠ��l�{�N(�����VJ�#�ێX=nrs���B	>|�
o7�g-"����A���;Cm�]Sߡb��|�i�<��[��3)�;��ЋSw�f����r0�n4��A��Y	��?{��� ��}�+�N�=$Xs[]�4�w%�����!K��wOb!�)p3K&�G�����!��ow}!��}���
�y�J��N������=����5���]��_P1;����T����c�K�f�Z�a�T�yvR���UfH�%������gk7BJ�DY�W���=eqp�7��4�GoD^��4<��,���˻�	]��ʽ����*e�q��P�K�n�q�ꮓ�j��V�=�,�yǗ�N�zŶJ�^�~�w�[(W^�CV��r��H��O[O'r�\K x�f�3�N��_D���<�]W[���P<J������DW�U�(��δM���q�^��}0C������[�7��y�֜�95��[�YMȅ�u��;�r({;47Ց猈�ǂp��k.�6�ܻ���9�VF���]T�ܷ�+zsr��>G�k�H�u������	M�6�[G�:�Tz�6�4n��<�l��+�j�r��uj����73�R絆��x����'7��ᗺ� !;�Z���;"�n��f]m]�U�حrn�Y�����}��|��k $�wċ|6���/JPz�=���D��Y��Wvs'V:؜�5�A�L��T7 ����n���R��;�dӸX�ݜa:��f��\�U���^�tt!��wv%����˃�MC�>�Vf��h8Rn7&�4SlRʸP0Cwp[ΛN�c��fVns��o\�0Zl�n����sv�p�q���rZ:>�����'�F�H�� �Jw[�I: ����9�R�7{�<�X�ׁ��/|w��Yk*�YJ�hB���!8��(��'�ff9�۷;߻T��e5��b5hPo>���K𪔩I�,�S"O�Ⳓs��IU{�:h�.gF`M/I����/����~�Q�S�>���|^�����xQ��^�ϗ�8�k�5��#�$P���Iy��8=`^�9ԧP�(ΰ�?%G��XL�U��U������S��ϟTZ�:�͓��}�|�IȔ��!�"p���-j�H��]��zrj��s�7�Ϙl�N����sJ.i��m�~��'�lA ���
�b�;�je�|���n9��Z׾ajn�;� X�C~q.yį\D�k��3�&pd֮pA �Hn��>��,�ȑ���z�	���Z��S��k�7Fzt>_8�#V��@�G+� ny�-ɻF���
�:�������ݚ�Z�a{e����<ք��fͺy:y���q��S[���]�=�gf��l�8؎�]����^M��`Wr&��_��G*軛�f��]V��`ٻ�ka�3z=${�WZ�vn۬Y4��e�:5S1�,f�̅,�����5���U}2�|��$T��ς	?V{}R�) ��� ���g�}�~-wRi�n*��-��F�a�G=�.�G�KHTw��H���%�r�N0_�ʖ���z���\�>M!�N�>ݭ��2"{>v[%5���o��"���Gw����C��lߺС�]��p������Lϻ%�W�W��4OQ#JbL}�B��`Q��>��(��u�kX�K�P�)yEǘ,c�j+�BH��fT�~��$c�e�d9�@���v�Gj0�bNZFi`�I��=��ZG��!F
S�1��+0}&���(�bE�G�2mpuY3�r��7����ﶜ|q���#k;�.��h�۩��DIإf�����
W���q�m��FA��+9�5��E�5���] ��\ů5Ѫ>���\�z����	�%���'������������Y�ԅ�����q^�b>��Z�*���D��c������#�ԩ���H���Ǌ*�I���#'a����[Tk���P��!�b/��￿�m�+ںc+�Ê��pb	��)��i|�V�"�d�|�=d���Q��7͗u��e�,Y�ln���ď�,8�E�у�#��$�{�3�R@��>��]�N���d�+�7�U�܃)�밑ҽL��z����w��	4��:�!��)�؅]w�Ys���C�a��Y�F�s'�$����"XIӫ}���ѼbnH��-�q���ܸIۗ@m۷�Z�6��-�J���UbYv�Z�|�I�D���\}��5"���B�	�\�.E�r>����ƒ�[��y#��K��|�q�u�D�Q)Y0�O�`3�y#��eL� A ��\L���
ԖP��ⷺ�\�-oY�c���oF��9���lR���7�&��2�&�v^,���);�������;H��cnE�A$�]=���>/|���Wk�����n�+����k�n�N��y�rtr�F�Mn̝�\Z��*c��L �E/��ݹ����a�&�je0��/Jķ��Z�g��v�r.�Ġ���K������L �:���H�!��)��j{�W��G&b޹��";!~����g�@$�#�06IRs�"�� ��{�K���Û;$����Z'�Ry�.����ؐ�p�}�a�K[��-.nn��Z��N{K/v�� #i�MJZ*YBJ�M[P�9�Ɇ��S�؄Tݝ�f�\z� 0��J^y��T%6�w���������<A/��@���1�����v0�\y��ӑÒ�	�l2�"1j��� x���Բ�_|����l8M��G#��B����^�>Z�Q9m��N-�1�����C�Hi�ϙ���x�Ud"8��[G֩�\��<M�� ����g-V��t�U�J��U$%�>-�.[��߄� 8�G}�~�m��]��%��mߒM�w��o	��<��-��>��=}|z�"+��	�੕��6��j�6�Hq�}��}~�����l>��RL�ϧ%9�7��ñ�c��=9�{o��	[�֞�>�݈n��A��䵽	��[�x�� 	�&�Ug�_h����ڣ4*<�:
��
+-�7s�3Cɔ���{��ڜ��������9��'v�}7�.=Q*��L$U�h]yQə��:B��1��.�o�������h�<�j�ܓ��#��@ �SI�!Ϸ�ǀj<@u4k���C9��.�S��ʶ�ai!W�͙-���-,���x�
ݦ�(n� 
��Ớ�n�\w$����{�.��>k]� ����XԱ��rF�ݔ�nl���bҥ.��$ja�C��m/z�Sl4��%���`�5�ܟp��Z�גt��k�"�N��d]�W��s���T誠�g#M8�K�m�A�3�,��!�����|����F��%���ɻ�{�=C�pFe��r}�Fճ¹�^;��{�H/9�ч���^��f��w*]b#���֗���s�lF�/�$����%m�z��d&�W��V]�M#k�9����eg'Q<�Ӱ��%�u��ґ�em��9����L�����䌢*Ki ]L�Wإ��T�лڎ�x=���'xF�n�x
}V}Oa���`k7��Ν�4_���x�Ep@�&�{���&�.� `e�k��b���l@���}�7�"���t�u�Ùj뚉��w���[�a�тv,�&3��d�U�VEr�A������=�zh���v�x���k}gދ�ŭ���c���F��}�q��n���_r���H�����v����IpaEAp}���]n��m�m��n3ӄ^�m�m`��m�ƶ싱nM Lګb{"v��m��ɝssnu�i�c�=�k�ݼ�ۃ[��ѵ��˃�9�ckMZ���
G�8ٻ{;���Rz�4�yvh����N�wg������|nv�T��Z�)�Ź^ѽ���;7F�E0X8���\��� ��utg����ٌ]�\��Mɓsϋ�l�:��
�1�=b۫���,�uu�sA���w!��pc��N�y�E�\
��ۛ���u����b�"�$+UX�⪘!C��f���ɞLוユɡ�ۊ��n����t�{�f���m��< ��X�v����<�g�o�T�۳W4�����{t�:��i�mom���ۇ�OY�1��m�����7a��f�^w��z�e��J��t�Z�ն�O�wnr���Fc˫˭���3u�y��<bz;;��K���g�m������zi�^�<��f�n���1Pp�{*S�g�%4+�����B-$�Ǹ9r��S��~]�2����X�*�=$\�����F�6��+�6ƴ��b�iD�dt*�Wpܷ;M#R*��p�%��ͧ�<�6�<�.�v���5V��e.]JEO6��w ��nfbt�ٹ�S�˃UnVl��8����J*d���2���2�����>�����y"Y]����<$}�1�ú�=p�o��wK}�
�zŁ7mUa��n�}Б�Ix��2�6'f�e+�
u|��Ⱥeť����m�L�G:�dba�D�.�U�&�ge*���r��X�@漒U���qT3��l렟vkT3��:Y.�lk�4l H�q��!�a�Y!�G=p�}����֔��0&����`��|r��zy��K2���ְs�v�Ŏ8�t�$
��ԋu��X��	M��	'7�d�w[��4Xa�wv��)�6f�"���i����0��Ϭ��b @K~�Z��uZ�[����Eji�$��sJP˞;����Gր�vy��a��+$C�>�;���&��6z�d�÷SM���Z^������ _��6��5TO&zF��-{�*�8�h/rO�=��I����%��0Dh�Dߣ�E�a�߫$V�D(�N&"UPU%e�IT�$�Qn����,�7s�.�&�)��B�"�'<�~Y���O@��(�@$��Fz���������&��.[��x�ɘ� ̯���Ӛ�E#��4�ޓ_�t��5ۃýT%A�{����Q���<ϙ��=ϥ�\�8�k|�ʋy&H�}/�u7ѥ�if���]U{&zb�Uc:����]vk�R۫T;(l�6�[）fbeی��I�l�g����A1�@����U'��|�$�o��^̤����Ox��Jj��s��g��Ć����:�GU��`�Z�����8�Ǿ�|�Ea]x;�56�5�M�n��4ܱ��,���q�ll�K���>]r+���R�}�Q�TT�\{��l ��T���H�̥�Q�9"���K�q��"m�<���$�j2� �n����
f|���z-��>�G��iG5�J����X-yףN�t�o`����@��/c�>�{���e�_�>����ѕ �D_�֠m����39t��U0/"3#º�lE�H5�y۔6ʜ��&����Z7�ꗳ����윶6,��K�������y�c���,�(�TI��,�+Q�.%XK�E6�Nr�͝�(�+�����%���8�iҵ�h�
�yU��_rN��D�;��S�a8�-��瀞H4:�޺Yf���S�qZ�ξ0���x�G0��P�B�����i�d#��}��F������������HJDq�i���J����ߟ���ͳ/@G1��=h��gm��\��z��ޣ�7+\s���K�+2�'hՍ.��m�!�Γ�s[���0n��f����Ngs֖Gu�|O��?��L�BGEl�J�5�$����r�^���MU�ԑ��*�Ic0��S�s]��K�]�9\�A��0� �Iآ�p�ԛq�y?k��W�Uo$B��q��^��#�Bg�z׽B�,t�=�����C���ߠ��jǟC�zU`%|��䒻$�ׁ����g���o�������������lh���E�*��Ŧ��]�_�a��%��聺�WϾ�1b���Dp ��_-��~�7Ҏ`$3��ysm�H[`��1��y�Z���d�|v&UQ�B.�i�v?���7U�A*IGk��,�PD��V���h,UO��=^f
���w��/�G ��������v��Bܶ���<[�x˳&eN�<�je����d�Ej]���p\:�b^��c�".��*��ȿ	*	�dߒ3k�o�~�)#HA��6ФE�Z�4�V��r8��-H�Άu�r��Q��Mn]�����RG*�J����|G��*Խm���Ԓ'ƣD`n*��s�aG���q���o�On/}-��S���#�U�N��\��Kx2�u�kѥi�?��߹Y�X
)��a\01X�sd�:[E#��]򒪞b�%��3 J�GF^�;q
&t!�9�N2��E��A~�z>�q3�64F��+@u���#�/�|�:�����
����O�Gl{oy���n������hj%}$��/7�MR���q�LQ+ܕ�IAަ<�R���N�j�i=�57J\]��{��N�����ȯ�V�����ϤY�k|)�k��v�� O9T�\U�.�o�� M�9�=�Ƙ�H'��pg�{��l�S��$�)�SF������x$�1'և8� 5�7�&�^��(�"� ��(f)�c%G�����v�{�>~;�q�&xf^���V5�[9�鲷����p9��j냫��9܄5ر⃇E��:tz���k���:��]y;q�9�=�aܜn�)��I�Knb���:�m�n{�a��1yW�YtO>Ϸ�<?X�5T��}�����Ź�S:H�"h(4A1nu&��9T'�v}��缷z�_9��BtOO�N�;��z,��Aw�,��s�-R鯾r���U�/i��5�W�o�
��3������q)���_Qp9��_imT�Ai�zv������;�{�����LP�"���=P����wz����E_��ZG҇|�I����(j�5ϱ�8��u�G��C������	�;s�8A��-:���*���Ngm��'$j�DL�95)�q�&��M�^5��IgX�Vl�^¨��ғe�Z����ڡ=�y�mͰ�2�d����Bk�|a�CW@��ߕ��uu��x�X��]n�,D%��Z�N%ʵ�3E�SZ߾��BϷ9r��η�RB�&g6w(��K�����	+8Ǹ8QB��4�ѝњ|�o���d.�$��;�cPM�|1k��V���1e�^ӊ@*q��&ef�J@{"�ĺN�D4�u�+k���f���.��)��=��n���n��u��WKfv�/�۳��DY��N�;�"�����΢�baK�!�<��m�"�tj�kY��	����p���f�^]����w��ت��k����Gt���`�����.qFF�-�}��L�B�3F^�5y�]�Y0��^��{���f߾-�,`@��u�i�����8�(Q�hldGlfZ�ۗɛ�7��ц�o�]���~�5QU��m�oaY;O����J:��jه2R��2�|�v���y�2,����0䦲���CX�d�L�Oj��̫��;�3�k+]�m�9x����s�����羆b-MQ�����Sn����Vu��)�sb�\�x�r�T����K�0�1�AǴ鲝De4A�oor����!7��Ȝ��,vf�	��X�P͌*��	ըX����MdB���Ɗ=j/+[�q��lS����v���%�h
�ېb��78 z�����&������6*��FN�oidFZ�e3OI���A���51���T�]bx ,7A�ϡ��0���Lƞ�M3�݂���2���*��}MwIď�>�]��pn,�ށj,�S+|�t����{y�nަp���5��{�fu�g*긳��Tgw�h��Vk���MpY�=��h;�7`�6'��x��L[���3����EDA����F�##h�!Hs�c��ƞo���Dsv�����sY�ʪ9�G��D[H����^}�|��9����qf���l��(Q��IkSuD���Y|w�1�	Џ:pw�J���L>{g�!�2��x�Z���T����[��1�H�S}��P�H���L=�F��&n�a�I�K����P��>S�٢��H��N�>>Ddz�ѥ�*Ӥ���|*6�t�1�'K�D�Ɨ�S�9���7P�~o�"k=�cbC'kA[B�ua�o��>v�z&�"�uE�2(Q;�O/�}@ �{<ς��1��s�Iq"��&{L��H���k�
u+3�T\���%�S��3���`Z)� #�"k!zR� N�q���!��a֪�U~J�q�X����8�G�w$�y�GPE�C��6�� ��]�#� ��Q9��]���H�����ت�r�r���7Z����/[�A�<��ܕW=���6v�v֌	�3ls���R����d��@[��r��=:<�C���eyZ�Qy:[�*�v������|a��: =��r�����6���#w~�����7�؂q7�O�#�:�q��ಪ��|ȿP���wn�p�H�x���hSW�~h�.���Mzۻ���1�\(�����2L{���s�+Ţ�(7$���|�]%z�U�h����
%T�W0QL�t�-m����u�h����'Q;��t
A0�Z�ć�y#��H��K�8��-w�|q��
���PN�$F�úU!%����ǖ�a~�4�sI��Z�w���6=̤�tj3���7#�@"��+(�
��C1	���,>賙�+d�N�s��<�0PN�|�ߔ#�Efy���fE��� �n�ه�u����2cz�J�c��5"��zD�$�rGٝ��R�v��Gvy��8��B>+\�:�}���DqjDh���_q+�'�T@��=��~5��������iw�M��H�w+3N��U9#�(�� ����0��t8mݨ�϶$�$g�U�#������JI�B;�����*�4z��~|s�C�Fb����"'A�(�p�a
��4j�&˚;䲱�R ���}�uM�|�m�A"��q}�E~�@]t>�h���H�m�֣4�湿�ܚ�g���gJG�׸��5�[����	FH�GѼ�����(�SF!�B��\��(E����.��Ԧ3���1u6S����)��Fn��h�����m�s���N�?���r܃�@��w��v��B˰r���6�R��j���"��QI<����n��B��q��r�;�n(b�9���9�T��Os�7��'<&
��'������Kgnc�͌�Ҁ����O�-�n|!���i��JY&�����72����LN�H��D �>�E�$W'�6��7O��ڑ:y��Z�|����e��;���{���V��ޮ�mn:�zn��0�'<mmq<�{uے�Ӫ�[q��!M��a�f�:��f�l� 獢��6y��=m��E,��V�'b��ѵ����G	��N:Oo�P5{�����}<��ŋ�x#c��xR���8�	��V0�m��L}�2�r:*�3��D��/��#��d(�DCq&�[E-okޙ�%���s{�i�pTQ���*�뀍j��Px`l�E]��{��V۝0"\�N憾�'N���>����$�zd�c��ҁ�0L"�A?e�m��coQvx���7Ȗ�ğb��Y^�3$v���P�q���|�I��j"-5��@=b^N땻CT��j�#�
�5^r�:�-��;�8Ќ��gvK|5~(�z�5v�c�J��ӹ�U����������W	��52�`ϳ�5�����*�������������A"}	Ę�����@�_eĿy���
�D�~9v3�qF���:ǧL�<<@]�o0GI`Ľ�/g*��Xq0-g�X4w֘M���nՠm��^����s@���>�L5G}�O:��? :�,�����{�|7.�#����u�b<�᳼/�VE)�0��N!N-�:&��W�Tټ��L��>�'}�Z�X�1�f|�n��V�!|lX}�xU��IC.���
�U�H�A��>���hӴD���T����*��`F"��JK\���A���B�H��Kz�AUN�}'ɠ����<���>�nBq&����`�y��n=��im:0РOĒ	�Bx��Q�ߙ�kq@_́�h�����5V������'����AM�j��ꕩG��0'-b���Ȟ�uԗܵ��)z=�"ǂ`�M_t�����FD���WC�=�����$���X�)0)UR�W���/�ؑ4D�C��ҎͶ}t��g����nm�T_�?��S��+����l�M�n��k��3$W�3�#����!2��ߥ���oF��C��F/!���G�i�L��K �x3S�lͭraudf�xj�Tm�Q�Kp�$�7��=�o/}�K��.�mi�]�V>�5x5^�x���5S*_y:�8�Vn�����w�5�ƢS���o���^qxQ���d����{&���{ױ\���W�@e�N���o��*�@l�8�����&>�)��r��+���dj�L���OMwc\��^���]�SՂED��>��N�3�0�hv�ъ[�3-�Ԉ5+R�޻��U�w{�;9䥦s�$�l�ޛjם5C�^t��T{N�KoI����'�{�'r+���S��Ͷ�}c�NqJS�
�xa��3QR�U�k�P���6C*$ܺ�ۮ�ڪ�+zOh==g�F���B�L\GI�Ս�[WE9�ͽ��zq�b��6+���3\����e�	+)�ÈMCj�ۋ�8�3��ꇎ{F�K.z]\j}%`ͳ�;r���!��l�M�n�]g�G�q.���k�E�3����cѱ�wcq+�<vx������`wѰ��+/��9���)zu��`ܙݶޖ�Ku���2�\����N� ����nx�]*8�=��n��v���� v�N*��1�ccm{�g�͓�n94�ۀ�����㧞�|@aN�;g��uݜc^{ �\k������ͧn���i���U��u���Lrn *���ixi�q8����]�N��pv��7B����;���Xs��ꞗ۞���\��:��O%�)����zt���Ѳ��8���Gd�喹�S�]71]���]���И7G5e����u����:3��U=c�9ˢ5uG����ùǮ�i��鼜�N��š�ڄ�i-�Iݭb�:�@�0\uaw-�*��<3�=ct�nx���KC�+:�9)k��zy�q�męI.'�,0�),t�j�H��c0sohv�Ь��wdb�1n�i�Mr�*�"Ewq����T��W7�:L*���ΧVQ5zWmN��0��Ƿ�Ӹ�{����8E�;w�G���BФ^I�V�|�c�Y�)�w*��i-���"<��'u/���v"��WE���X�x��r=���R��D�#�oWT<+E��Pw��Y�y�=֭WGWO�
�YA��U�F���
u��>���w��}�ǂ���=�Q/�J�x�7M��b�J�³SO;�l�y����A����p(�e��t��!�>7� ���)�2���0�oo���Z��˼#v�+����Iwl��J��:�nzg�y%�z�m��C����n��ۭ����uv-��r�����[h�n׭b�Z׷b�� ]S\)�d��ט:���Dl*RA8��7]�&�!3����}���W��rⲩ� S[)��t��؊��&�taM��a�h0ˈ^1Erk�s�ܜkT��v-�V��At�� �k�2/G�Q��K��&��-�zr�w�sؘmԿg��K`���.t-�����V�`��g/�X��i��qB%���Hb�k�Ϩ��=/�ƾ쒹
W49�Nwni��z?_g}P���>ԝ�~�¥�qT�ܝF�w�ھ�yz2�q>Mu>@z�	?6]���/�J�ͣ�E�f�������~=��+|�Ҹ�c�H=0�2�=X﬑�.N*��#%D�I�4��1{p&HN*�@_J9iz|�ObGי���4`Q9�>m���wꊇ�����Ҩ�EP�c��/s�;���9��D��������� nxa塤�Q�B|��4}J��L�����F-�;�"W��w� �D��Y������2F?i/D�p�m��mˍGiZ��軣d����?�Xm��۫��(��B�r!�����Js[����Af��Jp'��U]E�	�4�K��qphJ?RT�aX	�9dm8�KV��3Sɥi�{�y��׺S�r黊���n5庥��P��>��E�A?]�MB`л����A�#�Oڅ�]�~Y�r��K���W���{�-�%sH���w8-@�3���/ul��N̼��qA�\Q&I8�7e,Ȉr+¾Y��/J�#Z�91�/u�������0��ě�3f��v�-���N[XUJK}v�\���Hډp}u����/��wd��}�����%"����L��n�ϱ#փbaG��
pgؕR���\����ο���'�`G��A���:�~�,��IΑtjP�<��*���x�Z��"'����?L��*a���*A8	�n�7a7m�l�����sId6�8㝰����tF��>J^q `9���oI2Ƅ;O^�^.M������Q�y��N�{<�l���NJ�)�v@j���^ʤ�q93>�*c��U�����C��gO�����S��/����ȩS�)L����+t�H���KVx��u��V��̅r���I�H�X��br��LO۹LߐW�eI����+e8�>�FinR�M�+�y9�cuM���,}�Ë�+ԕm�>���	0�Q�$�!�}a�����5�J:QT�e�Ȅb�%��EZe�I˒<��MOr�wϓ�~�Mj]�N/-ê�%7�ah�����t�"n@��W{�peU�vb �����a�?t�$T��E�G����d\�U�(6���q
�E�kkyJ���T��̼����Fo ����>���؁�M
폩��x����
���^�"e�{��1��#�A�*��	�8"�\h�mgK㚓�ڐEg̶�e
;������|�J-̺�;��$Ӊ��0�\/Z]��R0+õDp�盛��,H�Q�GQ�H��ϳ8�w�$ � hiJ��ڈ��\b�/=2m���
%�Ƣ.�,��d	�RG��\���dΞ'������1��x�<�#5����&�����Aɍ/us֥:]�rk�B���K��8��zT��,ɬ���^���+�����p�*[�l9��㊽0�i�"��;���A��~؆��9�k�q5�=PE�9O���d��yC:���w9>t/�G�'��y��ѝu]K�S�ojv��ړ�x�C��'��P��J���n�)�>�r��'�6o��X�m�<�%oj��E�<7�$��A �%H% (���*"�eT�K:ӁUz��J��.,{N=W0y��J'ڰ*A$��,�E^�� ����CMNs�#����(�7�>Ԯ+1@��\`}�#���������B3�n=bw�z����^��Ǳ�Y�=��QD9����Ϯ[씈3#�!�F�h>�i��n�W`'B���F�t���i�-���٧���7Du�-�z��n7m���B1�-��Z�����l[K������֡�u�-�犎��W� an����ע�/�Q��J�P,���� �5�1��E9dv��7�۰?K��m��87&�����HE�ᶢ6�I����	�$�P�v�\ bn�}�M�>o{2|~�7��H�Q��F����sw�'g|�Y�����.�eג���?�� },��:�u)����:S�{�t~em����0��\��B����p&�)�5A�'5�H�a��sZz�����e��3��<����O��#��c���������BO��H��U�VQ��Nb)�<�B+�8����a3����!�6�䦷�5�\�-�^��J`������G���*q�[
04b"s5��U�F���=��$h����G�G�i�]��s<����fa��#!"�Pp�"p�:'Y�5K�8*Y���=dC��ȒI=���ð��n��C���mג5p1�k���႔M�.ՙ��g:�x3��I�+��~V@(�^�+c���9���j�,]	v�z��ʼ8Z̾���������~�����E6T�%jd���}ד��tY�����p��V��y�ݯP�[��(���5�v��vj��o(�M���ڷ��� ����U����V�,��8�T����S�F퓻����=��tǵ�cS�oj�5�89�re8�w�.��6",��ϵF�7,SK`�f^�g5z1���g��N��r������d����aa�Eogl#-H��ޱ*l;��{���͖��[��\(���Y����1����*2+���[��Sji��q��yB:y���fm��ҍ�ۇ�+xO9�ʽo+{!8n���Y�fE�s�m/o{rߌ���y���sh�2^UZ�ˌ@t�	us�s�N��b�g��rU䈎�W]CA�b�9/s>D��[��y4<ͺ�X`Өj�9k�kh��A[��(R:~�v+*S����S{���;�����-D2�7]�ktAVa���F�Ҡ.��N��_a�[[w�����h
�7�Wtvf�o\��X�0�5��!V!3�E����J��)��ֻI��+�����'fW`�n$(�.��j�ə��)���ꠧ5�����Q8�)�Y�cJ�(.T����=.�!\`�ܱ7sw�|��k>�u۸�����sk:+�Fݬ��qhir�3qI6S�Z'���U!]��;��"�GH�����Z�a�Ja�d6�Zz7��(�;�tFȚz�һH�Jա������+l�b�E��y�S��u��֯��I܊����'ZL�,4�7Q/Е�b�+ѹ�2�n"MrG�ιK���}"塛�m�ة�A��y�ns�nn���.�#u�Gѥl�n=puS����6���t�H�H�x�_��T��0b���.�����7��3���a�ˈ���j���l��b �"�{C�/���H�)���$+��.����v�i>�:,�f`�ύ��Pw,�K�1��M^A'N$��]�G��ڬ�ߤ�����S�y�$RM#���@tg[6����C�88���q>�7t�/�\�I7�Utg���
*��v �9e��B�[b�O��j7��'1#6�|~w��䏤ݮ��kE�d���������F"'���eH9p�Ǌ&z�0>�NH����B��*k��X��<��{�LBr��_?������EǦ�^�X��/V9���H��m�6�z{���W�<p�5�=�n��1:ۈЁ����u9m=m,x��k��f@�ut��D��I�H
�r���U�6���d+�E�����!T֍��6ɪ\�ɬ�zCV�ҵ���<�5t�(u�Z���H�}q3]�#4������=֜��g!	N�7�]<�z�=�}�6�x�ܞ�	Uz�խ���z�g���(�ߦ�p�佂>@���m��l-�$����?H�ح�^�|fN6�n%��Ђ����N�e��g��-��_�rFm.�{�M�#V6��0�Q9���D�"<���'��q�]�P�� 3�����T�>6�+�ނ*��Q,W$E-�<���N1�pjΔ~����/D�(@&�6K	�����q�B�A� �7П�f�+��wЁ�Hܥq�޹�"��DC�w��bZ��|#�,k|���':��eB"l1@&	��[�y�4&�sGܖ]7�ƆĐ~9�#�X5#�Xe�p�2E�_�;X�d�{ѭC.y���y�`Z�DMd�.t8� ��f�?�W^I���{/��(���{ḛ�yW��61�j��܊31d��m��K>A�g�_J9*��r��Y/�,����:N���A�zi��y�c�s��a�SnY\,[���)GjR*��7�v��6���|�.������πL�$5仩�B;:���'&��.&�V
�q�	�^j�h�U_57�߭׽�4G#�`��Ǿb�D���Ԕ�Q^=���g<r�?4�~S+T�~�Sm��r�DK��f�9("^�����K���ג3�u�6[��N�ѵѨ��t���5�}{����s^Ľ�"k�2D�z�Ր��m��9�r��[}ic">U`�'*4��=��m�څ��,�=��l�$�;ڞ�6o�-6�7з�¡�b*�d#����2}io[q{��	 G<@0�5?�*����(!�r�.��-�~�;~��4�<O)�ۣ�Z���@�����u���ǎ����tq	��Ćzp�E+�U���n�f)�e�dpk��y�Whcvr���^z��`��)�	^4�dFbq�ɯ�1�a���J��{�#�*�A��E�d��j Ye#�f���t��=���7Ϝ���2����w+��nN�W���;	\.��xU����?;C~�H$ͣq#��W&���ɹz�7��s��Y+r�k�(��,�j���7���5�N`�fpFsE���^n�fcї�D	�bhD&ܷ�W#�3|�]7ϰ����Se�P�Q>�W+�z����n/m�X&"}�s{�S�~�n1@`�2��į����L��#R���;��ΞҔ���ݥ=0��;�LtL��k�]�ؠrR=�y�ʏ�q9;AqTsЌ���R[עfx��%�;k�?o�D��U)b���h���I�Gܵ�Q;���~l���i�=��\�),Q1���X�V���B�6�p���A�����M� ���	�{�C�l.�(�k�d�XG�8�֪�Gk�H�s�y 5�@w�}���D������W�>$2#�Z�ݜ�a@�t��z�ad-9�+^)�ynY莂p��ؾ�8�{�g�#4�""�5���}�7�~�0��z��{nYd3�r�/��ޕ�e�:���+�|���*wp�Y�vΑ����ϭ��Դ�EQ�B3ILA��u�l���㮫�{`�a��<��}*SZ~�g|��-��OVzon��g��m��qnI�>�d�:;�>G�޻Ev�,"�>��>��?2���O%�
�۞Q�oL��m�Vm�u��OW;f��V�
m-�Csn�jB�M������Z��fw�-Lg���D��`�A������#ۂ�1�{5)۳�����~_'{R7){o�zEA��X����P�Q�.�8R3�Gi\¬)x�I�{��a�5y����9�>8�U��#v���q�����Kb�^A��ԑ{�]�f*S|��I�T�����GR��`���ƚ���sj���/�ZFjݓ�(���� ;חh��؃�3��k�cG��ϸIM_��Q��ŉX�5dX��hU�_C1.�K*{hخ�U�DV�腇��{���:�����*_D�}˽�Ob������mV��N�ڱ��xhGfa[�7Lq�}��u��6��.C�q��vS4:���Y�����c�w6
P*��*����Gj��8��Li�U���E}�?o@E%�{
������0�nSdn�X^� @��� ����=���_�3(W ��L��j�v��\lg\��{to]2x���*��A�O��ɾ�ӭ���P����2��U���9=�vH���AX�T�a�k��.��͙v�<Q=���t�&��+k��`؜��H���Ԥ���ń��5�	�=���׃[�U�/9+.�����c�g[gu=7/\4��[���7V�`��ݳ-rv�js��8�0݌糞ޕ�R:.�V�����������g��!�Fy׃�%BѰ��>�0���ѹ6��v��9K��V7!#��Ō�nn��棵�����r<贞n��Wo=�q��g��\P���u��6:.��3���<�=r�]�;�wTX�sgٙ�i޵Y�&Y᱂�[��T\gn8I���tWg�IS�(��m��1�n�������x捷*덹��r:�;sưr.��wB�͵����؁4��2��ybd,x� o�h�l/ny�ĝƪ�i������\��n��3xݤVwn�����7"�n�)��tH4�6��`�r�:<���T�X����n	�%I��q���[�Ƚ���R��:��jn�dy�!�q�OW�	9��^�8�	��c[N��<n�]�Evb	O��"�E�v�^M]����V�K�cM�Ac�Kfr�[۔�|ws��qd�����&���_m���nd&}�u�|�k{y�ռ�-Wi�EʛI̹��/r�y��Uw��t��Fv�j�d[�b=�k�H�gJ��j��^�y�%���TJ��S0��� F�i
�j��E�n���!f���@��wI�+5�U�|�QȖq�ػ���X,�t�����}�L�����q���Z�Z;&f�%�YR֩�Ŏl۱�-C�i��j��C�u�Q�3��$n�T@۩�7��,�ל�� A�KzX��z��l���S�q�Eg:؄d��@Ƿqu�+��cuu�w^���-9ʹn�f�Y�1�V�T̿���Ȧ�0b�$UG!*��(�qx�p�m�n9��'m�<��]i��i��v��EW��Bp`���nx���f8�&�N�D1�X3��Ѻ��<�>,�\�@�ӗ?xƠx�����E�K��\l#e;��Te�'2&��C�pw�Kn�#3��A��9��� o&����紜A��@T�l���uΏ�Ʒ;�1n�I�A��~n�m �b����L�#�H�غ3@�s:"��8e�{�TM�]H �Au%����Q9��#�#���m���g8�䛁�ž�|�H%̑��K�9M���w���mV �K$e�j��"���H��R�d���w��`�?���$S��g���9*�y���xZD��L|�5��&�d|������;���:��7:�eF�zt���̃u�����5�8�J�]".;�"l��9)s �@V��g�Y���梦+�����W�߭'J��^C�a��y� �[�,[�>�5�׷�u��E��m���@n�B�I1u��:�J�����>���'�\�����|�I�Y�!�r�g�ɞĮ��@+VbTc��ʬ�=@�GW�"�_QA� G�2G���W���F��&~�*o�xL�}��G�8�x�� +���^G��a�����a��'�{�^bFc�@�����I1�	wg}
�vԉ���7u>��r)���ZN�*j	m�A�Z+Z��Ҙ�3*�B����!}h�&����ϻ%�֟}�U`�c~ďR������g<����Pd���R[F�G�,�U���&f�N)���@y����]�W)�@�� =����]�/��ʲ�m���$�	���6څm�u"gU�ȩ}bfL��M���Y*�Xl4g���c�w�z�lw��'
�[����d�
&�G���Z�tڄ"E��}��ߒ�Hި�J�DU���E��]��D�5U�{:�D��^�-���gԕo6}�j!��$Ǳ�\Q�>jH��߸��ۏhU��ﹷ���9��,�d�­`y�.}��'aD��s\n�BP��Z�y�l�9��Ԯ�L�=:����ں��8�V˞ܝ��qZ��rc��b��a��F�G�u�e�.ZWG��s�gn9��+u����#�'H����O?w\�h�ܕ'<�76�f	E=6��3�����0�~4��z!I�������-�7;ٸ�u�����v����H��/� $����QD7���ց5�+cӗ�U����t|��^^���R��5�7X�2+M�(TZ`��zy��#�>k���I�{���L�{�,�+OX���U��Tb��������&��̫�f�w�G�.�>�xH�^�̵׫ab��Afy#�� Z�'���� ޱ�D��Su�a �}]jd�U�"|�t��9��1���t����5r�մ��-��u���+����8�\�^��2�}��9ܗ ��$㩄}o�������id��o6�}�s�o�%Ak�	>]І���ioK�!��Z��-�K�mػ/b���8�ԌI�,q����nh��H��wahQ9��6A3i�"�X�'�l�/7j��+�|�z��̐�V`�Ul�g��ai�߼H�WNfRbLb@L=�ڌ	��h�گ�ʰ�2��A^���]�q�H�~$N�~���c����?���9�:!�iy�c�:�!�r�Y8E6�m_^����>�e�l�b��>d������>j��;��y�J��{9H*H ���GB��U^�J~dщԸx�F������p$��E��oj�J���h�u�}kW!���Q;�D1b���>�!�t�L�8��n�#��{D�4Dm�]$��]UFܥ؂I9����L�v�Zo�q<Lgp��;�vMNzr�}����}9l/�N���8R��	�1>�7t����2h����0]Wyk�&�a��6g:}��M�m%�'GqH�(�1�}C��e���i�����h9X��_lC]��&�&Q��]񼀺+�余�� �<�@�2y��
N-b����Ӵ���'}q��ٹ$^�h����)��ض�͐Mk��gы�{X�㳖A��n�],��;�uV�a�:�ۭ�i�b�ۥ[�����:ۯ�.ܛ�nt�u�~��k���f�s;���CU��e�e�I$v~R�~�M�O���t����"�8N(n�8��#�8r�p]Yɜ�J�9��z�z1�硿n���,I���$�M�U�n���U���Q`ļ�d�=�"�H�;�O\�*V4/�o)#t�S0Q��ጒ"���� �7ש��mO�Ř��3��n�R����š�?N���"�N��1u��'7��)s�-�У��f.��&��9ߡ4��
?�2P�� @ "0���rjy@��ͻ7�F�9Vz�p2�,�Z�x��xf����T>��73�����|OE⃰P`��$f��>h֥]Gѝ�I���R�ڑ��$ق@|������Q�${\���~��"t����$�;H4�!%UR�"eQ�*��z՚F��-7�Bgv��k4����l▐��ב��H� �x�P�R����N����E�Mw�n��76*����i�f+=��^8�� ��Zh�k4�<z�z�;�7���{�gC����
�&�c��;�F�*�������$rke%=�(ܲ9^^\�;4+P�5#�n/�����ԅ�Yp5�7a������ꚨ%��GO-Έ�3�'��I�*P �r�ڠ��˜%��V��3��g����+MpN/��˚#���=I,g���|ƶ��̈ey�ۧy�q����0�Nww����W�b�-�nwl)[C\�Jξ��'�Q����W�o�<�{����)ƛ>��W�3��v�Y�!<}n8˻�$s���

��m�EZQ�;-�Ar��g��{u�^�c��N�ݯ׸T��V@��}6(��9���4�v���c�����o��f�=��S�[�[sԓ�/�e��t��ǧz��\l-����#Y��\1f�T�h�H��쾘D��x��q��(���ٱQ%9��yyk%���=�_d��Xn9wZ�e^Z�wͭt��V�Q�1s��FZ���;�p\�����9L�,�j�`�r�s|.���j�Sq�ft�@�1��:�a듆Xs1W3Wj���Y�Oh���ۂJ�9�9ɓ�@�jV�ޜ��@�aNؼ��;�.w�Ngl9.�d�fZ�[T�9��Ÿ6��5�{������t3a��B[��[�U�s.lsj�/*[�<L��nd�v�k,�f��U��":��'lf��d��&E;nĬW��()��&A��!����þ��e�5#�X���T�Uk�m�l����f��ؓ���i����V�N��N�,.��~�����u8�o�����Ϣ(��f�|Tu�}�d\�w�Y|�@8�Gjz���	9�R}x���|�8HNy)�|�v�=��q>�)���9l�S=5bxƃ�|C�:���ی��	>���Hd]�؁[3W,P��;s�^�)H@��wꉲ��U��LHX" ޺����N��Y�{휎�*)^;ø���`��s�e���-ш��o� �����F`E �����ߛ㳮�`�9��`T�k/(cX( ��⬑n}���Wt��t�̦!�F�Ǐ����6kaT�w��D'*��-�ə ��i����C�(%4/����R|qmȐI{A����e˭{���7�^��CX���'c�a���5 ы���bV�|DL�A؈�M��"�*������ӗ�\uj�X��������W������EI�]���ӹ�-s�U۱`=�����'fz��Լ��U��=S��7GoNH�k��_��>�삆(�dQ�[�����5{��	�u��4ӵTp�Z�Zq�P�gC�pbٗ΁�I���'�#�:e�4r7ࠀK��zz���$�
�0�7W�n�-D?�&����|�q����~�"��q�K'�(2o'���	��v1qD��!���r�g���ǰ�r��v��f�Z־��8�RMB��;��~����y⢷��)���й��_�;::>��L�l�v��@컼x="�Q�>����[02&�'�Xo�2��=��n;�X/��ԯ8�`6	����p�J�ڑ���D}%�6#=��1�[Y�����=p/�޽}�I��#��"�j�T�B?M���UI�Q��w�^b%����+P

�2�;U�\)q��Y���Z��yi�h�1f6���"*�y����w���v�;����\�l�JNr�|+ �+״ h!hn.�C��>@��|(�O�0?�l��q�\ia��q�!>q�Kh_�Y�4�R�1�I�|�jຸ�SPW���{������j6�؇��r�K�=�jN<o��=��?�;\n��"��p�r��+�V5�m���M��Ꟶ�Q�"q���b7���A�fE,�o*��:Ph!�.u��O.1�y�d8�����F��-!�z,s�ovE����"����?!��[�ˍUJ����: gծ.剋�v#��&�Dd2�bIP��dNV�^����)�"G�}٣b!k$�.�� �9ג{�����#�5J*\I�֩)P4�S��f��72���/��o.諝��F႗�f��/� ��3�V�+��p���z�hy�=n�"H�M�~;������8n!]�]�@�$�U0������]
ɾ	�MP��H����9)w��RG��y*?G�d :2��M^��q}��k$#�ܶ(�nF
��C�+�Y�0es=�۱n�f��z4Vv�okp	��u���y�t�ݲ���l����ʱ�zM�^�<us�)n����Eͣ���&�M��4�8�q�Tbg�=�X���1�Q97�(�;���q�S�&/��	Vó�2 �M��z\�$�]͆������~���+M�ˠ�D������i�Aӯg��9mR�u��D�;���^�t�1'�M�s�3q�E��N��c~�,a�ɘ�}b/��E&�ìž��G˷��j<Q�<�#�8,����m�������'�^���o�"�;�rsr��j�1v��'���Mkޓf��|���G�k��*@|�!��6�e�8����©��m��������(F'���n���q%�W�pI4�#��	7���@$�W������]R<.�.���rD��'���m�ns�߁�1��A�Пlo�l�#�Q���2�]�qd`�bS�$?E�w�̻H�� �����oDKm�~ؾk�ρ���OS;����K1o�r�U�����hϲ����G������g�ޖ�y��NM�a<tr2���Y��ֳМ]�������Ma��ST<�t=eC95��w�$Ifx��6��F F��T{}7�~ߡ��mq�X����rؙmp�)L��.Ғg_E�4{>�͑�_1{g��5g{s�+ey�@]��	"��������/�E��|_D��;������-Db ur��)oV��Xht��GQ�Ru��+=-@�H��L���b��3䉪���T ���r@��9��-É�1>��V����M�u�%�'P�uIT,�A8��EyA�ӹ\�޲_u#����\D{�$��,�S����$�����Cl2�sѷh G�f�Gx��s���,��9�VGzW{�@q1<sF��T������F�x~�� ��Q����%UQ������p�>��f��}��7�:�t�Ǧ�:oG�9�2�1�	)NK}��ТI c��lqm��b�a�m�1��3nl����F�z���:Wf�`������߆Ơͻ����S`u�l9��͎�g��8X���٥��')������|!�":�-�sӝ�7�s�pm��V�͍,PI���e����_����~��?տ����}�D?!�N={�;�����μ�mn���to�����v��/���WO����χ�{_����8�������zw�=u�����3m����ח��~<���v?ߧ;?.��-g��lh���Y�7'�oY�_O�?O���7�n���|���9������~O��4����}�����f�36ߏ��;g���-�o�{:����ܝ �����Y�}�q⛩l����<7��[����������۷M�&��:x�����������|�s�����r�~OW�硅�m��t�a�B"��B"&�$CE�X�D��-��ɢ��ȶ�&�-d""i��Me�D�����F�,�-�-dBȈ�5��5�YY�!e�2-���,��-me���M�k&��ɭ��DB ��-dșY"�Y�l�h�!d"�,Dȶ���Me�-��-���e�Z؈��Yd"�&��k-�a,�Y���L��L�Y���,D�me��X���[D�Ȉ�YZɭ��DMe���,�"�#E��d��Y2�F�E���"�ɢi�DZ�e�ZdBɢk"-�e�"�mk,��Y",�ȶDMmE�"ɢX�dX�D֙d�me��d"�5��M��5�[h��"Ŗ�,E��-�e�M��,E���e�ֶ����-�&�4�!d�"�,�E���,��&�[l�,�X�����E�����Bk4MY4X�,�[,�!e�m������Z&��L���h�"�",Zk&D�,��5�k,,�-k,��[Y2-�Ykh�Y2ɬ�Md"4Y��E�2ɢYD�L���!�E��#E�L�i��l�Y�h�ɴX�l�e�"i��d[,�L��-5�Z�4MhMm[,�E�E�,�4[E�țM2,�ȶ��[E������[Dk-�e��me�B#YdYY4L��M,��"�!�X�E��D,���M5�Me�4Me�F�e��E�bȋL�i��dYE���ɢ,���Me�e�Bɢ�&�"[DE�Ae�MYb!e�-�œZ�mme�DE�[E���,�4E����YYdZв�h���B"�k,E�Z-�Qme���""�X�Y���YD",�&�Yh���&�YZȖB-5�4K,�,���[E��YdMh��"�-�"�(��Yh�hE�DY��DZ"Ȉ���Y"ȖZ,�ȢȚ�kE��Z-e�dVMh�k"%�YQe�Z�,�ZȊ$��e��YE�,�k(���Z-�e��Qm�E��K"&�d�k-"-�Y��E4�D�V�ȋMl�",����Z�DYdZ%�K-Ցi�[E�Z(��-DK-d��h��EkYDYDD��ki�E�&��,�$Vj-e��Ћ-�k)��-�Q-,��$E��%��h�H���E��Q&�VQEe��%�(��-d�-e�,��-5K	�Ed��X��Ċ�E�Q"Mi��$E��-dD�Y"�dVZ-e�"DL�L�YY��Z"Y$Q&դK$VQE5�%���"�"�,�������[I��(��,��D��e��"��+$S(�K%��dE�(ֲ���kE�B+)jjV�^\�nQZ�)�VJ����T���Ԧ��-���EQ"��iiZU)J$��UJUj�j�Z��%Ej�R"���+T�R�UeI-$�R��ER�Uj��Z���֩*��R�-*ʩEj�jV�eJ��,�ֵU
K��թ[SREV��%-B��DYe����K(��DYZ�+H��,���������h�)�Qh��K-�-��D�eeeQD�H�(�ZڲY��jŭ�ed�kYEb�bEe%��X�Z,�5bD�V(Ւ(�tゲ�
-b����A,�X�Yh�+VQEeb���,���d�b��H��H�$ڊ�2�b�bD��-d�Ŏ4K5m��YYX���+-+�(�H��\p�+-6Z�ĊŢYE�M��+-ee,�QYD�e
�kb�%�XLVղ��1b�E2�Ċ��&ȓ++H���!&�YF����Eb�d�,��$K����2Y"LH��",P��V(�Ykie�ɖ��&,�D�Ed�+-�-
%�%�Y�d�Y"�BƊYB�2%�D�E�ME��X�X��+DK(��"D�Vj-d��bmX���D�md�h�k$HK,,�Y!Y!&��f��Yh�"ȱb�Yh�(�Y�"[Z-5��B2+-�"�e�DkK���E��4H�H�Yee�m�KVZ&�D��D�̈��d��Ee�4�ekD�",�Z,,���mY"�Z-d։d�k,�H�֋me�Y���"YdFYhZȋZ&�,�&"�Z%��(��mh�D,�5�D�Y5�VLDMdYY4E�i�k-�,��&�,�H��YDZȋ,�Y5D�Y�Yh�&��2���,VMd�Z-e���D�D�Y",�-����DE�D�e�D�d-4B�"YMi��tv��K7.N7�-�G/���~.ǫ�?w�z:sc3m�pb��}g��gv�����7���������#�����)�{�g|9߻������}^�/�_ճ�?�������1�6�������_��������՝��<���{;o��������_c�}?tu[��i�4:z���^���z��u��|�����m�fm��ӻ��f�;�=�������<o˼Q����|�����=ǿ˷,6�k��m�3m�����c�_�e�.3��Y���rכ��{�.�xw8c���=|m�ͷS���ѽ)qˏ����r��l�[#Y���>o��:�d�Ɨ��B4a����8 ��<Ce"�׉�ɸ;����6��_���_�e����y>;l��Q�����}[�� ���y����g����>`����7{=�/</��&�V�|
>��������G��~s�����:���ff����{B��h��{��};l��pnN�p��=7���>ξ��o^?����p�z�G��|�.�-��8/�����&�w�3ƛ��=?��{4[M����_����o�v��<n����u>E���?o��o=�fm��S��=��8q�V�����{�q�����;>���+��xݼ�����k�}\r�<u�v����z��p��}O,=���o��l�ͷ������L}��v-�����f�۟���s���:o�Ǯ�ϛ�w������?矷��Ѻ�?�a���3��rE8P�9:d