BZh91AY&SYXE�3TI߀rxc����߰����`�� }��@)@�!@   $��Q�}�         (   ��>�A@P �B����ǀ }z@X_U�٣n���X�����wl�ۗ+�z���=�\� 	��nwz��=:�ۂ�*���A��qOZ���
 =� a�[�ׅ5����o<P$����Cx{׉{b� QRS�l�b^�vi�:�k��<��z5[�� (�=�ëw�A��ި�;��{e4hzмsqӣ���m�6�x[د;:7gv���8�C������P  6W����4/�h�����p�94b�Ih�Aû�)M��$u��
rіA�� �Pz��^L��P�qN�Ol���;�tK�G�T�P�T�q@�z=�C�7B�2ѡ�                   O�R���&�4M��D�U!�0     O�*�Bm*  �  �   ���	�*�@�L� 	�CFCLS�2 �P�&4�A���	�a1�`T�D=A2�S	�<�=4�~�B2z��zj��{���G����������;_lf�b'�����i�ftfͶ�6���?�a��ɵ��������_�<�����6��M��bfΛ��{:U^��Ѷ�l�[9#ū;�M��o�g{���?g�������������:|{�lo����e��)�Y�����M�X�[6���æy緎�>�����8ux�|>?���O��O����)�p���o)�4��9��T�I�L���_&�#�mf����{U�d��
s�**�D`6��f�k�UJ[�]ӭw�n,�/����%�F��0;��:R�_+�skoKC![��j�e.Гrem��V�U7�2�˱�V�[��ʢ�J�ɺuH��D`ɝ�fL���ܵa/����d�AO3��4���!����e��	t(u�����[j]�H�X���Q]�gγ6e��&�Be��zm۵�Rő��i+!H��peμ�X����!60�:H�v`�O�⯅ѧ}\-�
��ƨ�7���7�2��M^sY\�[�Y&��7mLd�,��/J���7h����{��J��仜0-ou��[6���`��)�l��]>�-��)ovJ�X�<{qԙ5�t�2����4�aV���!S(�!�B�E��qd����Pv
�'���cT5���n���6�S�cvD��v�8��r�ۇ�m�△WF1V��v2�3Eڧ���.��9����Nj�:��!u��(m�\�0�nE�0=sT�&��l��3.��eZ�h�]ӴOt����4�MF��W]2+{-P����g'i���o,����������(E�l�"��n�ŭ�vkѕ&��8�v��/R�inћ�Qw�u�m��*k�Btd���4�T�9dfC14e�he<^6MZ�%�](���j�XO10��s.��Y{(��&��0a�)7��t���*�˶ ����yonAW+*ٖu�ʊTE�j ��r�lm����i8
�6̖�(�E�*�Y�'�=�����`�F��~T�nm��ث ��'��Y�����
���,��>��M�Dvpf0�+V�0�˒�hȖ����6���6JnH�n��f�zp�Lf*���F$7�Kem�&n�,�����8^푴�`���~�,�i��T���J�8Ba�fD9	[T�����9(@w�H3�2#�e9vj�
lG�^aV4�2�-l6֭�f�F��g����̫�-I��X�E0�����ku�)��%��:0 ��N� ]9e�8zv�%NhP�$��y����Kѐ�M�_0SM��T�X�ǊT�6Zf^�&�Ȱ��ͱ]�M��wv4����+)[��"�eXԻ��-a�I@K�	��Y��mۺ����˛]-�Tnh5v.�/J��F]�I��7Un��l�t�Ņ���˼�K9.·z�� w��f'ش��pޝ{C$�)H���;�iT���滭.a�!������5��[W%cQ#f�`az/v$�������9J�ܘ����Ͱ�U�*6t=��d�vj��n�)�e�ʳ*e*�p·��� u�}�&�ܶ`Hk�,�C��ۧ)��Qfd�1ZX�-آ����#U���īѪ�ï()l�{B�pS�)�b\U�o]	��A�76c�a���<�,-�u�j�S�F޽oz�tk(��8m�
�V�Z���r��ڪ:�7Maw5Z��t���o!�mD3��^�o݌�th��6b�o.���77N��GF��u��"��˓/�#脎�e1,ߍ�����Q6�a��vP{�^X	:Xȭn�隘n���^��ƴ\��Y[� &ݵX��ҳV��u�v�a���63]�������d̹`	q����V���Ʊ��B���4ḥL�Z��X�8��Ǖfd'v�����X���hQ��%�7��K@Ѻ�n�w�φQ�j
ˆ��H�b���PŨ�tj�"BU=���&R��T�/�)Y.i�ܫx&R?0ʫbQF�JVFcd �i�͋����ָ�ʲ�I��t4����2 ���x<���d�W�̝#;�Or��� ���Օr2�y$aZ6ku�n��̡}���'q������r��꽩T�qXI�5f�C$�`!zb��8�C ��πR�h��Fѭ���u4
�0�}k(�PWe���JΓ@�U�v`ܩ�ù�v�ik�Z*�l�KN�&���bt�s�)�8$2!	�J����
���a6U�7�����R��WIV؆n�Y��N�Ȟ*ᨍ�⢀�C�U�O�r^��X��R��1n�&�8fd����/��1��,[�3,["9î�r��a|�\�5t
����%�&%(�7l]�g�ۺǧ3�#;3�!!��;C�$c�T�.��:�ͱO�����`�«nhm2�����O}���l�(�I���;Ѫ����@< w�ֆ�{;vY��1J��9��d���P�7*^ԙt�H��o0�vLcF�rXbZ���.�sFMX�s�I���Jܛ�m��̵�]���������8;�:��r,/Fd\��)�)�Q3T������3b`�h���z�q�j�v�� 4��K�Ż!vT�� if5s+ �uwsGi�M`���!��Hk�%$ī���N��g���YUp�X����TQ�u�yT��C&��aO3�#O���en �j���iL��ؙ��v�}����믎��־~��>�u������o����s�y����}��<��+��H����Bس�o/?S�1���F��ɭK35�}�V!r��Ka���ir��N18�(��NȔ-���:q�/�(V��8�[=�����-�>kq[Wa0��	�l��|��Xx��m�v���^�#c.�у�<�q�x�}u���ɷ-�.��\֎��n(��\�^�+���cu��Ng��f����}]��]��=�7��X4{��%�ӗ+������J�k�_O���l�2�O`:S�{9��&�!��������}��9˒�r��\�Om��sb͒%����a�[d�|�u�n��CP�Y��u�٤��<y�^��N��������9wj�)�{Rl���m�)��������c�؎=�NI�I�H�q��<W��/}n}�(��e�;65�[�ֺj��.���;��f�U,Q�	1m�����:Ʋ��ptn2s�F��.g=kzz��jݸ�l�¼������qFA�ō�����kr�(t��@�c/	��$+��{Z�����^x�n�`���,#[Kvs�-nα�����w4�:tn���v��mq�]`�zU2�����,���9��ԝ�9������c���ۍ&)ڌXG���$��Xx�j���/r2�^��g��	a��C�B���1v�ZL�����^�N���퇞y��]�Z���]��cm�upuԛۘۚ89|2A��-'c��m2���<���]�i[-�8=& �ksշ����U�ps&خnD՞���н�ֱn�m��)7����b�QL�G����ؒ�n=����pmVN{I;n�tlq;n@�#���z�dv�2�W���i٫���ܢ�%�ێ,'xi%���l��-n����˻9=k+�m<h1s�m�Wf��DQ3t������gX9�Ŵ�� �1�Q��s&��\�' �ی�=h��rx}[�7)Ihq�������`z����v�\l��k�v�A���F4��V6��ݻl�g[���h�b�:2m�l��<��)�Ѱl�����;=���*ޚ|�#㓘M%�/�v�p/�f49�"-�:�)�.��Y�c���s��wj"Ө��mӦ]���&�u2��گ\���=�#q���F�o`�v�3�x�z'�6m�n�{5g=�����x�wYyO]v�t�.#d����g��6�"Ҍ�Bp�ֽ&V�������	�E�w;�J�[��ۇ�����6��WOq���uG\q�0r��E��!]C']�w/j�F3�x{\q�G��)�M�뎸}�ܛ�G\�Oo\���b뗥�OZ�s�Z�ƍ�CA���%��Y�:�ێ�ݱ�ʻ���{��O�;t�ͨ
f�ڈ�Qi@����M���5ٺ6� ��N9�ؗ�}�@��9�f�����yk�n��ݛ�N�/m� �κm�ڠ��+����n���Ŋ�7G[��ū����<� �2n�q�c�ܢ����8�k\���\ns��l�A�l�s���8,����v�Y���kn��k���F���,��f�3�Ճ]v�b웳�U\�)x�g��xN�&�u��7�o�v��79g3�v��\�'k���V�Z���q��)WGU�(烮87�s��|�\m���݁0C���6�v���f^j#�u�r���JO ]Y��]�ېmɞ'n�������/k��(��AvLmK����;(#;u�Kc0��G�s���t��s���:�S��F�{C���on�[u;_v��Eb�s���jy�y�i����m��c����]>s>����7�]i캹��<c<:�z8�5y��mvh�`�]�vӃ��uF;��m��u�u�V��i�k�����>����w�װ���������߯��<���ϳ?Wό��E���~_���!��'���̙�����+����gz�toOHʥ,m^�[�[������*q�E�*���fw-�6�%���jr"��|�2iiz�1[�C�A�p�2αZ�1W��Z�״�hɩk�ݥ�d�6Q\�C�3:T�G��nn��C�CldNb������DL��1�l���)�]B<��#EI�e]�qj�V��{���:�o�E��,�:�{���rF�ާ~"�d�կ'2�d���u������[=��F�nn���;s.�����\���Y	�Y��o{j�n����;+��*�za6�K�v_`��9כ'kY����엫���38ZF���2�T�W�i�k��$�z���)S��Jڏ���iܮ���n�a�W2��@��v�EH4J=�v�GZ+5u�"���q�����J��i���{�2� �Ĳf�;�/;��+�S�+J@�:'7jf��)�k&ň8�a�0a��K��hkz�1���]*i�]>�*����aX���Sz��.�%ydC�&�:o�{��vm]<E�N����k��qw��W>�Ξ��ܽ�J��*,&�S�k�BJMgu���:8HƯ��\X�l�㶱>1MXlK<�t�wv8�'l��i��ٍ}�ؒ�SǙ�o[���"�(�n��lY��=�e�Q��ihh� �@�ۙW�-���NoE���Z�e\��EW]\	s9V�< اW�6���ǵȷ\��{z�=r�]]�@R��Kw ����]�8v�!��Y�t3��;n��\)��-�jB7�U�G`_9�pU�b`��0d�30n��Y���Y�Lv��fcBfғ�"�,kv��9rԂJ��׻���:������9	��b�۲�3g�h�� �c@�Ig%~�+��4%EiIzo6V�z�n�#vK����������۹)O:�
��EبHʳ�5�gB� ��B�p��V1��^�Ì��#��j��g5��t�WcY�1˞p�X�ѽ�����(N	Me�l�13��ǝ���)[�3q,�.3�����PP�#}F����=��.���l�+E�lT��]�� �l��u=�y�oWo��B��B�etm(��ݖ��z�oybӳ�b��x�wz����P
隋�O8��S��e��}ڦ������,��ڴ�)��)s���!� \�X�y�ެ�d��5�^��O��4(�1�U�
y�-n���][�.�h@�IKl<�E�`�δ���%�C6ܡ�n[��hn�Ѭ��#�v��%,��R�h��*��0�'z���n�%V����v���uڨ�Nu(	[�,N�G4���5ǐ�l��e0�Q�>�0\R�V�dG��tI�n�&�n2�7�P���PUnV.�@.f(�p��Մ��a��׷Z����[�᭰�e[�mB�bߺ�Czt��ŷ�&��t�ۖ$S"yS��O�l��^����7$BT�kl����[Qm�:�Y�Љy�l�ZڌY^u�%᫸�]@�a���s��W[�>�Y�V�7V[���ɉ��x�ɜ:=��{%�M{J�I�����G#�v���V��+�Шó�'t�y���=�ř+��u�\]�����|	!}�� N_m���T�+�y[}���1�*gMr���iS�#�ahk���Wm ���Sةv��v���fB�dV	z,��Bd�2l�Z�x�;;lJ5��Ѻg@���6 ;3J�ı�{�p;��J{39���o�%)n^v���=쳳����F�M���fnq�p>�]vs������w��=��L���M�	��z��K�����h�7�WQ#fhu}�Hں|&��J���6μ���kضVsT�32�ݎ�GY�oWF�f�j�����N|���5M��z����i�%
�m>��P ��Q֙ע���vG��.B���XЇ�n%��MH��f����*S]pVE�+xŏI�R���n�-�^��MJ��S��i=ù�~�!z����ً��F�AAJ�m ���Y�̗W��+=F�l�3�/�k����u���GҥGO��Q99ڼUbW�2���[n���7d�8���7E��'&+řNe�ƯE��U�;�J��ѱ��cF�cзtG�b���B�iw�)f���&g[�@��
��!7�n�Ya�G�NU.���=����Iز�r2�Vv� �]������X'��#P�xi6t)z�rd����YR[���dt)c�E'�2�Cխ���]��f�pdu��gV��ҷ;7�Xlc�}�<�h"g3m�C/�EAWHn���5��}�V/��Q,����h7�j��=a�D*��%�[�]���V��4��yJ����*>���]��5�H���׫�tuY�x��C`cvjown.{�c�����c��.nC/�yS�*!gE�ݶp��
���� Ł�][��1.{�n�0k/yS�e6�3V^����VTr:;[���B�z&S[���{��gW%�/��̬�D<��v㈝u;VJvwc�}nT�W7���ZN�X|sǎ�<;��ǟ::��oq��ώ`͖�m+��������_�~�Y�>��	����8�|m�+w������U�t����Ӆ�v�������ڎv�ڪ!fށu��z�f���������>>�^�UȐr���n�!�K�����Mw\Z%ݞ"�;���gA�;i��l�n7mX�к��</�m:����X����$���a�;�K��q��Ŋ"Y��R�Zl֛��:�sʀ�q�g�ݝ���;�I�&��8�O8���c��p�H5ƶ�"�۶��햰�b�.8��s�����`����=v7�66��	��lJm�<����t�Wv�
s`��4G �۴'n���u�Ğ"�"Z�zx�,I�!ۃ4���m�nn61��ڮ#�ϧ��d6���^h�u��H��u�&#	�������	ڹ@L�.�MA����9��U�h�⵴ql�ӗ��SNݸU�3#���û͸m��cd֖�2�	�-��I�c[���-��{:^���Μ0��T�]�U�>�9�/k�ow��(���`mpV�'V
��dw(��+�E�����ij��p:����n7�N,|G��$���c.7O�]�Չ֢�(�e��,�U�U�"q�f!96��F�o�ws��]��V���Q�ݛ�An���!���Z��n��[Z�{����DSEN.Q۝����5գ0%�27m�l��s�g�Ass�s����ƺ[���t���S&{e�;gq�8� ຎx�>��v0ʹ�i)��Ȩ˵��C㧢���6���K�]�����%��+�8���/N��K,BK��Y�?b��**�i�֚^7#�����hZ�7�u�~����W_�R��Ӧ�����M��:�1`X�O��`(	�=�Q�~��[i�=ʻR�dgv�^���;��w؏b�/	S�}ڴMq�k9�EN0̏E��p�ֻ�煬���"�}��0�L+�,W��(H�,����#�x��w"MczX�X�x�>4��	��Tr9HQ@�IK�C*<��)�,�Wt�[EӘQ!�}�Ʈ0ҿ>�p���7�Jߴ�S�"�m_�zgk����ي�@Ĝ�b�	8-	D5K���v�ܶ�ފl�z\�&1���x�Y�>�,0���6���a�|0���+4��̪�X�Im��u�����ێ��{���)��vٟ#e-Y��Cv������(߫.��*U~�����jU�w��{���T�m���%����!y���t�`�F��j��H��,�M@510�����:K�J'+C�`��h`W�G�� �̶�#R`�Z��f�.i`�֦N��Q���$Ģ�6k~lQ~����]����
�H��g1D-��>>��/����"� n�����PJ�c؜�`~T+���tW�*���f�wg�>��G��w���ℵ�
�X9U�OI�,99!� �eu���y�qW9��d���=��<PV��UMEX�X�4XG�B��p���,�[b���wh�X�Rj��"Ž��r�A �Zm����#����+����g���kJaT�W��fI�߁�_�|G��/D���0����w��\���3{_L�,""�����,�"��R�ug�W�<��;M��<$&??}��|����n����U�6��I�)MWb���Idr�ǦRIQS� ��6�yTܡ�坢�kY|̢Zh٥7pm���J���W���|5����?
E��~�xa֑�:p�*�?�x:vk����VYPu�M�f�ި!v�v�69n	ujR"QЫ������_s}�,D���!�˃�6~�	7w9?x4�{gv�׷7iܽ:Ɓ�y�='ֻ����^=1X'P���e^'����s��t������!�Ǽ~�d��`,���.�	oe�e�]����L�pĢ�Q���
kX�2�;_2�.d�64(�X)yU��!���֜#H˕~����=�yj���°{������z�Y��L�z�0��=Z���	+�lm��kHu]J��!X��+m�lW��\7x���C䏼k�ɛ�����h��z�ua����P�,�0�gⱈ��o��V)� j�z0WC#�5<�J��}��x�����:^̣�t����AWL� �{�#���5z�}�q{�L�&�~�c}��$�c�Ġ�넰F%���N�X��9��j���Î�4�yx��q��:�zA�������k}7)�g�$��(slc[��~���O>�a�Ӵ"�XX�".f7b�C +��өR1F
0(��Ң�p�tY;��>������L�,8]y{^}�SJg�o~��|���%�o�(��S	���70��F��+t��4���8M�pݲ���Eq��z���@>�B��d)�X��7�z�ݹ���h��~�'��gd��OR��l7�K�hWJ�Qd��ܤ���
�
�{#���.+�T�Q�K^,^��j�E�B��KZ){�>9��2і���Tk�7ߓݦ"IX+iYFKM)2Y�-�̧�>���P7�$Y�7BT�
�� j��]o̅��/�~{��؄|p��o�Ф��2�.��&��jͭ޳g���aJ=����v��l����qh�F70��,>�ү<w���rI΁�>��ԑЕmsz-U�iǝ��-�����7�P*]���#�Awc7{oM��>W�Zs+����P��+|��,�@�g�|w��9��id��i���ut넃mnvC��Y����)�[.�{��������m[`p+ܺ���7ө��o^��ɷ�&�׻��Т�u�kNQǣMӱ6։���jX����:�-�2��}�����w�q�̗og)�ˇ���Y�Nm�G1+�-�E�W{������^E�Ď�������f4(���J��́�^��$��MTL�S����ԕ�f�7%����\\�//,V��+q�י-Jq|D��B�`�8(ؼ�a�[3���9@�)B��^+��&�b���PT�,�M�b��Je�%�f>[�)���9aB����A���i�K"v��So!�b��#h��#�gu1<��6�9DB���fۙ����z�j��D�:��+p��Ut'q'{qo\a�r�����pim�ΦZw�@�-�X�.R�x�ή�xF[�W9wJ�cj��`�1�)I?��T��Z)�؊��Q>B@��ď<q���Ӂ����.x���:u��ٸ�V���a͏�&9��s&�ӛo=9�#qo���K�t��7�8;����w��ͳ����N�m��랝�>tch�qGCЦ��"1��Q�Ӯ��n���ٝ{s�ڳռ���μp�g�.;����v��py�\�8fz�9���]��4���Ǘ]�N�����&t㍫����K5��4G�հ�����=hL�x"<&׃>��~���|�Hf�O3G~�;���>�3ϊ^j�5��P���}g~5}��e�S�1D�\f仹��5iP���nf�c����ɺp�m�z�3Ş-��寛{ܞ��RQ��1KJ�`�7=;9���M�y�)����.��-*~��^��{���П E���!xHw��ͳ�����<y��\MOޯO<��v���X�<w�t��pីp���{�����h�>@��`H�&W��x��;SQ����q��ۉ��}y��<�:����Ì���^�l����[9��6���(�y��WGej`�6������'����O*���y�M]^�0�)�jܻP�&^��n�V#Esݍ�O�����f�;n�n�;ĭz<]]�1�g<\�^�yӝ��<��8��qe�h���,҉�Q�o�4���.:8�I�v?c��z��]׎���{[]8�&�g�<=����9�G�׷�x��N��8��oV��W�#����<O�#�~��@E��獸�����7nmN����
sӆsm�n,z��۟Nzq�v�����<������IX0a}�����	�fQ�&׼p�cˇ�q73��7Kg�<�ݦ��Lc8��W�V���[S�+ac�m�v�#4&���{d��φ��a{l0��H������H�y�����9��s��6�ܝ�g�=IúF͸�n���t�:.�[^v�=y�eo8���ͬ᝽/�f��l�p�e;��x�I�Y�n�8��'�Wn<��\x-ŽX�k��=���öq��Í��z��Ϟ��\v�՜[y�Î��sV�^��eo3w�3p�u�8�8��t��T���QVݮ���Ma%�q��v���z����k���g=x�Ǉ��]����<��㍫y���N3�<�����Tg����2��}�i����5���wyC���͸r�~���U����
�Y�n�N8��Q�ڕ��ԅIA-�����5�x>�Ïx����U��ۛ�~7Ke��ZE� A#qx`�/�����I f�3��q�<w睕�X�k�3�]N��O^���\nx�B��ޟ˷}��*W�>���	(����V�=��D*e�?��yg}'DĹ��e柂����A ���$��6 ��-z["׽綑��H�i��ASY�`��2o)&�?_}͛�R��J�Z���ws���A�v����{���+5���p�P1e����!*SD�e�/�6i*���:ٌ�Y�5�Ng�g)���Cл�A��Y�n��c�#((�,����!�3��$�>)��u��RycD�����R_L/��V+��D
zV�R�[�B�.O�+F����&9z'��=�7OM� f��c�=������!�;)ա�{g��]�Z˷D�Ю���~�uc\��ڸ�8C���1O&b�vO��M��F=R�c�f��-ᕨ�Ѐ\y��t����tEU�R��ߝ8ܙ��I��&yR:�=�$<(��v�����ኮ�͡�(Af�7_I�	T���!t�BK�Rs>'�ШQ��M�<e��X����<�:����*)a�ٙ����<���C��|+��ً�x����	�qb�D}a} �L}4��L0s1v�B�{����k�F�w#�Y�2y�����-�3s�3)d��+�ӊ���C��U��H�cﳥ�)j���J����y{�P:6�pD����W�.�G�����4ʌZ:)-�(�jLTv���H���'�љ��{�?c�exL6��{�����gB��Q��L�����AI��}Wf�����t��$Θ����^hy]��:D��s'���Mn��P�U-G[å����/��UxS���6~CJ��"y��:�+�g�W9$��\�W��A����n�z$�]u����طc���`�b��b���Ûn>胨H�c��P����>(O6q+�4Ê�|C�6�� ���&Z�>t}����ߢ�	}���o7]����b=��U[Q�~�G���~$��b+u;5R���ij)7�g�����[�~�g�<S�^�)fCs��
;����
��|3���r����{�*k<�0�Q��V��36��4�zԮ~1�1����x���n�CK/���<�>wJ~��<B?�'��q��drA��
���T6�7E=����5<�r���?7�0��+Gn�]�p� ��n����=i˜�Q�G����1f��U��e�%o��)�@���^���7�!r���j\�uiy��ߠ��ٻlb;:�+�-�㉘j�U�޹�=JZ���]ni���]˖��ʤl0(6�ӝ#NV�+���r,�f�3�������V�$eҦ��Nł�iӼ�-����q�YH�)��"�]�Z��loPܯw2E{��߻N{�]6���9��*�Ii�Ǯֶݸ]���[h��I]��8��۶q�&�K���8�S��{W��n^��n|<��Ԅ��
�>�p�۳ׂ�9�א���Z����e+�g#��0	��l���ژN`6�k�;g�Y-x�n�mvȶ[zv�:�ťF�ܷ���v��;����b2q�ضۡ���G+P��q��XL�3ݔ;7m������Q�uPpV�dۢ9܆x��i���9K�x��a�u�\K���7��y�&]�w7A�Α;A�о˹��Q7<��x�ko�͞^������vy8�b���� �j;�㧞x��3P���<v�W��-��$��/��m�n��4��l\����	�]��
$��s��{��L���R���?7ϻ�vmb����5��^����Xu�G[����U܊Z��8iW�ݏ��J.V_�_>˩n�R��7�s��;�;лNI�ޜR�q�z�/��Y����V�Z���MZ�ͬ��ˈ:՟�������J��l�]U�ً���6�U��:��}��y��ݥ�L(=kU�&t�	�/h(��F�͚�Av����2�-�k����SdS�]��I�ǲs+�z��zmƏ�#��Udb��ǋ��kn�����ÞR�8Źx3ۄ��W\M�0��y�ι�h����v�?��-�;\��%Q��3K��y�n\Ъ�R������P�{-� �n=�`E`���RHE�������3���@��������|@�G���u�
soR2s��,�}0�[��D<�#l�>m�� !;��!�[z\A<Q1)�u����/7b0T(Q"��e�r۹��������o�YmI<\j���9ru�4�
�=[p�����!�z2�z����	�����SX�i2¶�7y��O���O���[�a]�;�q� ��(|�O}��;E�^���9���wb9�������,(�+u��_����8xY��\`��<ܑ���i.��F�f;s�[œ� 1m�\Y�r���4���lM�y��&�T�&��جٚ��Q�`J<
��?c��8Hd���q�)F>�NbW���DX�Q<U���hEW��0k[<��D|�C8m��Q<Q�!%�͝(��8���0|�#���Ҥ��Y�̘��בBK⚜<&����VQ��;U�ze]����ut8EYC�q4G����'�o<�����K���S��,ȼ���W�1��ݙ�0]	b����U�G���jT�υ��nɔ���s��8���'->��v��Q�l���r��t&�q�FEI�#��I�����OTY_l3�3���K�����Z�74�RP� Q�7K=C���*���e7�������#'�lD,�����:Yc�9���l�[?<h�����(�|���j���T	�Rb�໊��wލ����۸ش�g��=�E'��6ٝɄ��*�<8]��C�F��n�!�"���UEsߝN1���bβ1����i�9�$H*����Y�ju�gl�a�m�^_��������n{�'�ziu7�ۿ�ohI�D�UM��8�_l2o9`L��7b2ۤ������Uv��U(�5V?ٓIw�eØ��!�U���`�P�(8,8�x�Y_uh�IҚ=�3�+�]pwy^�������O��?B��	�Si���	P��r�~@\��
���i+�B<�L�
�s[�l�'��1��&�f~��Yli1�?%)b���s�M�Z
G�b��=�L�簐�J�����}#j��v}oɸ��U�E%
�)9	�����#z�??�ju�ݪ0��5�j>
*�d�R��T�s�vb��F-���mA�,������5Cv�T�$���V4�x딩Q)e�������j�KCƯy��|�<H�{�� ���0��X���vy|ρ����:Q�"|c	L�U&�dM	���<���٣{����]�Rςu_so��2�ݨ�$gé��=�f�x1;u�]�����W�S8U�r�
e�ͣ���u��׏�\$t�U¨y#8��Mt+�+����� ��;^͓SH�ɉ����TMK*}ݗ������8�h�e)"-Ǽ>+�23�B!xB/<xn$�;�� ��:U W�j��j��%�H��/��ؚ�t�,,�7>�q�e]|Tt7w�`x+!4`�sS=���S��}8η{?�{&����n|�g�x�ow�㫉v��9:�6�鈷�����v����mW�����ﺮvG��q�m�c�;�f���Gk#ښ�3U�y��.wo]�(�Z��D��m�E�,�=O[�e�/u��ԍ�z���Hm�$_�\�3kyO���9+��=/}|5��[���7��!J���/��i��?ksM疡U�h#h+'8U[�Wc=M�3�L�\/`'�G|!����/$�Žy�~+� ��9ژ�,P��ʬޟ�VO�:��X����>��k-�mB���"�K���{��W`f�w!a;[G����E��]%�sZ� ��E��ʽ�3���j|���G""*���!�aA�˘��Hx�3^+�kg�n��3�٭�R4m���D[���G��ii�l���,���SL�8�$��w�oR?�>�,.��K��+`��S�_*u��x}��<�-&�����R��O�(�}���{�j(>�n��+&i��`��B�W9�����_���x�D�2���thf�MY����qaq]�ҳͩn�}t�r��P=y��]��R&|vY�|�^��}`�*M��	^D�}o�+�����v$ٛY�@^��g@�wSloz��w3yg��ks�g;�u����vp$9�$�­S�ߋn��%��x|0�[�6����I0N
�7����usl�o�����0��WC��Cyi}�ˡy�jS���$
�h�i-�J��p�]��t�ؑ��.�M^ʖ~�1telL�Q̴N̩P�Th>뱟lٰM;�lp�d:|��ͻ1ر�d�f9��7�չy�k6�&���s�η�
ȸT��K�z���P�\�{L<�wu"���3��
5�*CR�qh��b��J##LD$)��9ܸԆ�V���&���"n�Fƈ��w�#YP�H8�1N����ʹ3p|��:�|�˛����F�9i��0=bWd;{��l]�.���nA��Y�0D�K9b������V�=G���z�IV�^3�f]�3�_]�(f7B�����ȝ��+v��l�#��7���k,��������21����_td����#�k	s�����vىjuЉȆ8��T����͆u)��c<z�[���K�Ժ�ߛ�ǈq}�i��`���� ����au�9�3�*�'���w�[c�f|rkr���BV�����rƶ�.M�,�5Ĉ+*�Qx|�6��*Z%��kۡ]���kO�?,}5�>��M�)�#��%8S�Q�)S�9U!���.�_b�(�r��uG� �*�#�n���3�l����4V 
��8��z�C
�=G��],�(���;3����d�͚���Sm������)�*b��~���s�u�O���|�"i��nQ4k/�.��味LM�]Ǔ���]�:�ku���<.�[�n��2[�Y:��:6�V����+��K�_7���V:���,����oi��8)%lm��@0��K��_�&yY�>���V��'��Y�(��G�?6b��G�o-^Of �c`DNx%Ŵ`������F����Q�#���o�{����"��m�S%n2��� EP��}&�;���,Ȕ�CAU�7Q�f�RߠҾ\�~�;�G�%W[Eϴ>̓ܩ�]F]&*�P�2���Ld�d�k���G�G"��6o@.�{�Ҝ�T�& ����ql�=��|!�s{�w��uu��K�ͯ�����85%T���)r�4��w#��J��<{�nI�œ%}͜*�덽�(�U�_u�5*<�&h�d��zޥP��r�;̫;3��Uh٫]��#��	�(�Q~B���d����7- iR�}�t,4�Kq��k��ሇU�6~����Џ���Y�(��"69�)a#q0��E'%@0��f꾝X%,�[=����4qo�w��(Ƴ^'�AV݉"������ ��V5�q��S�K����vF���Pg���7���`��i�.����+�AV+x�H�F��+�'�e��-bI�a�B�!�#����9�'p	ʇ1$j
�U�
��LA�=�����B���(���2'�{��ܭY��΂�U_6M���	�\z��f�Wkg��Y��r�;����4oXo���ɒ�eC0��iG�9'��v����� mp���#.��"���!�D��%.�s����r�ۆ^J+����3�~�⾱�˺�:4�\�YK���"�;t!�շnFyx��z0:ծ�eN�~��p1����ԩT�anv�Եk)ѿA�2�p�z�$��QN���[uM���x�)��
��	*��`�Ȉ\�c����0�$�F��G�,�G��=��U�t)������ѷ)"�w�[��q�Ϥ�Й��ߤT���rGP��N'F=�FPo]��a4s[��%�2g���~�rb�����s姧>�/� h���D���^w�i���2�4b��͘k�Ԗs[|	}���bѳ�(����l�6݈��=�1��[>
XO�F�0ա�K�!>n���U���>NT�zeP*�*e�ZdYS6�����������hX����k��6���/*��Û2Ww��g]C��ɋ�3�a*�E2뗪�Eܰ}�g<^aR�r���U^+�7p DH?pND�,D�k�R��;�bMOx�����*G��9qV����ny�݈��dH��P��e"�e(D+h)��̫�����G��i������=�3�#r����=X��8^Z<`��y#��l��縴�&JU�I��#/6pnn�oP+�7��D�t��+�*���EF79�j�Z��~��p�Tq. E�w6uo��}i�L>�4�m9�ѵvԵ(�͘u�����,�ن5_s 
Z�h�W��|:G�4���[4��`.����7}	Q5�Ҳ�"��m��}|�o�����&
� �Z��/PΗ#��9������E-[z1���hś��T�uZ�Y(8{�3�
p*���s�%7Y�]���Iuw�z̶���~>���W�[�3=��ջ���|�_f������JĜ�/^��i�>��e���LRF~s���]�=z.FwyfOmj"�-�˝�h�R$��m�R|���ht���z���r�'�ӧ
����K9�}ֲ�eFϭ.��9)�q�k��������Hd�]F�����Y�pnX9��%��3*{�uf*糏W�%Xʒ����Z�{Lw�|�MM�yp&�4FV7,a��:�Dg�%I�u�a����O�P˲����Wu�����q����)��ٗ^�.xވ;&h6�8v���f�۱�����K6ɀ�NzW=�]��=��H��Gxܙ�r�ۧ�>�G,���'�c�k��Z�sԧ�N蘃��Zn#��j�َ�pv���{��σ����|:��)�񫛎�/\^;h.����8=Q�c]e��۝�y�sVl;<��l�^�+zX��I�k����NV�UQ� ����b*!P��=��vN|�M��=�O��on��Z�uvj^i�6��uXϠմlvd6@n�������V���uȹ7��z��v��rd�O	�E�bY���ι����=��K������m��8��Ywn��x�3@*�Y@l���[�njy�ua��Z`���=���ʨ��=��s�@�C��Kk��H�	�]���ؼ_飅�ۍs����Q{)f��튣�m@-Kb[����_^bݦ�Nvm�����4η�CX�f�2��.9���w�Ŝ��,��K��{1���݌�v���Jt���o��UH��V��˚��ؒ'h����
śU�T0騩����*%ԣ��l���Ͱ#˶M/n:0v���Ѹ����װ=mӀ�b=����z[�v�R�a��2[;���{=�1�T㍮5�����q-���"���~�n�v��\���#��G|l�v�ϸIݶ{����*������al(�<��{��L��&7����|���z�5���tb��l��z�&�ߛ��/����Gc�+!9w:�~^�us���u�+�D���Η�"j[1��$���z��J���?:u�.Z�7�ht�y�5L9X|�=/6*��۴0[��Z��
({RU���>�=�Mj<���*�����B��I���*f�S��{�$�Gn�t��#���u<<�Ym	d����U�m��l��B�N�w��/��tm�]���l#������0X�J���'��N��U���٫ƣQ��u��7 �����R���� ��&!��>�fފ`ก=��[8�stlAχf�tMZY��Ti�f��}�~��g<5�Jm#G����swm��|MJ
;�N3���y�6a'���˺�؈*I�!c��t<A���U����o�nF�<o��G�5�-?��\=��ο�V�XV=�byl��;���YWM�M�j����~_LY�&���xa�����Z��o��L2X�5,�T)�2K�I�����VSR�D3��!�¬��Xx�A/���9����������>|`�6~Y�ۈs���".�AH)�'�k]US��iqI䞷!����{(�ZNs����*��֫2'y[���r1�j�Ud@���9PW�s���Q`x�i�t���^����յ�ݽ�:�q�⮈�س�*
�!�*cy_Y>�����<�I��1AKjϙ$���hi\j�]���#&]A���vĤ�� ~q~�[��UЀfq����U�O�k�̤�_t8����D=C�u{)��9�H]�e1�.D�]ܷ�1�@�;X�c�j�a�X��R����F�ӑҍ�w�f�f嵿��w��)b~�I
Ψ�Md�ev���>�}_�`����8LCo-�k3�����ǂf���iNѭ#{5�n�ml��"��}��d��uH�V�r0i���]K����Q"�R�8알�=�犵�gO��LeBqR9(��A����1"sܪVl�������Sܴ�g�Bݯ?H�65���%\J��6+Z`�%FL�U�|=�Q�k�|!��k�1��2ma�F���rBl�_|�4���U|���k�Q*��P���'9�� M�"��ggf-��H�Ԥ�&�f��Sfw�.�� 1���c��܇���gZx����k��C��uk���$A������]/�U�<g�t���LX���1sX��+욟��N�G�w����Fa�E�d�o.�ܸ)F�}�b�JOηJ��f����OEi���F�+��h�)���$λ谽����c"�]��O�b�@7__��r� ��A�&�/�bk�>�W��놧���@*ӂ�+S�ԇ=7\�Qck#m܁�8��i�JQ(�i��cc�у�%N9��Q8km͝�2t=��n�룠�:����j���76�P[����u�Z��^��<$H�lR m��L%G�*!5h�lw#�� i�c�x���[��0G1m�a�Ӭ�#��w?=����?>���	�=�:o�Cc�ϜH���˷Z[��;�q`;���H��Y�p�b��p�/V��Ò�ýrgB��Q`/mw�:���u�q�'S�</IU|�h��Bs��#e�Ă�QY��X;�,���f(���((-�(���X�;2EC��\!���RU�~ڭ=O:�j��M;Js�@^��}ʳ���5R|
3�6#P~�]*N�x�����2���h�Xʣj=EnG�_sg��Mz=���eD��>�зW�[3�5�$Y�Xw�L����_9#"��1��U�=�'{��[���7ڮ�!�
1Ohf�k&�w2��us�r��\Z�7�^u��c�n�
�s�8;�:�������z��R��d��������Z_,�.b%x}�����G��m"��X�Yj�hKR�*N�%��qw VP��v��Й��:	��r>�N�U�㹷G&oKPG�n�"�Z�}��2VZ�f+���p>5wԅϒ�ӧ;�G�тe�.��x�=�$�]��z�~�[;o�����b����e��2�J��F���!:���vV��ʹ'�*f��^��5�9�%Vv�[�r4y4�\�7'���<��]�*n|���{E����\onqdǴ2�Fcb�^ŁR(_���:�e<Q��r�9��nr9�α��F��vp�.��.s�Y��P��z2����z�@��T5�캛�4FR�{��<&��2Rip��A鵹Y¥��4�Z�����?���bN�xi֞]̭�d�z�u�n��f����%���B��ԅh����V�PXab% w@R��#뤗�U�_�yG����B�������0&�z�����E�q�IEp���8ںK6VL�����<�&��Z�j!O�A^�C�CM�� um�0ڞ7Q����!q��߼}��,���W�҅�?r����r/c瑘�ؚ�w�#-S-۱W��皥�lW1��S&2����kW.�jЈc>�c��ʣ���<G ϼ����Y���rS!�
R��R�74K�"0�$~��RQ�>��DMv���By^��=��T�յm��qx����&'<��E.3�B1}'��M����J�X}&����G:s]8ݍ������}q�-}h��p��p܎{u0��g6&�(��ˍ�䇧�.�I�Xn]r���^۷j�3�9��`;tO(��^Z66�s���(�J�:L�2bEi�����PW�u�-��(g��W;J���y���$��Wf"P�Ne8�VP�t̗���>���k�R�՛��'HS�c�@W#,Þ����Ļ����$珀ϖj}�������p�_c�2��'w����DĂhQB�&��5�X�`O؍�G� ��U=�=�28w����h�V�N�v�r��#��_���\�q�����*w�.z�#
��8�.ݵ��3���H�ʜ[Xߩ���}�5���Ǿ����)�Ǐ�܆����� ��.�P�M���W|� "9iS��ڮ,��jv�E[$�2���V,�2���=��@��,��D}�=���^⑇����sLD�+��&��r�>��w�mU����%���U�T�er���fn��s7z=J���"�b�r\	" �V��-ɣ3���V�� �+�t��"�������
4�WpY"G�f�y��w�3�o�%j�RV�UF��wM���z��'�|�����xT�����c�uR�R��z�xA�����I�M��
+��-�O�?#��vܦ6m��N4�į\���Ec�b�T�|ɕ� �=!�$�[�bȹ�U(�!\H�b��sLI#�v/a�Y��E�|�RȜs�ˠ��_���&�~78������M�~
����Ƈ��^@*�V�D:��q&�oݶ��<|>3�U�|4��(tNx�^����M���_-��D��.ݺ�r�lH��ص6�y� ˄�#W+�k�u��Ǝ��q�s��bC�n�jt<�c�nE-b�V�s���q�Fg<�Y�����s���������B���h[�h���h0�jQ�{JgZs_\�i��3�J����R���%V��L���n�fw���ؚ���������`�xb�U��W�O��S^õe!ƀ���P���)���!�hq
EM/M�sՌ���T�e#uQX��D�1#��]��+����9��; ������$�L��{������I�_\�ڑ��=,Sl\$�	D7ȁ�xa�[�k� �J�h*~ L|�܆��3����a9d�����UÝ�7�޳ҷUd� ��6a���88G�U"�޴��է`��xW֦�PU�.�hz�q��� ��ό	�T-L�{���|�o��/
�F�EG\�oM����˸�ؙ�
'�������ݶsQnq�ܛ����<�v!�.ꤜ"�H 
�}kg���GV�W��
L���}ہ2dZ<G���>kIo�K�jQ��Uj���Wk�(&a�狅}��k�x|z��6!�ܴi�^�8GT?�2D{�+�,p�z���Cr�B��p�1/xv,/���fw�߻S+3�w�'B���7����JW�Ot�XL�440�b5khyRjd9������)�Y�@
����IX��Ed*+��)E#B�k�D���Shg/y��`�}�<�qV�H@��݄\�.��{�a��3������*����k0���@>�G�	�z�B����ʊ�+P��4M���d�r �ꗴc� ꇿk��9ґ��^-���2T��ۊq���t��*�ٝ�.G�]d�k�c��Yr�m��\�.Ȼ]��Q�Vd�[:���\���W-o۾]/ީ�	���(
�^f�����C��g����X��yj�����w�U���X�����@<g�1��f>��h���fvw��`���kګ!
.D����]�ۥ�}޷�Ϙ��U��`޻4�S��À�ʚ����r�y|7���Z�_JgGc�<o3*	��viC������&�n�P)ͣ5|�~�nW+V���I"n�H�JJ�yWp���N���G�v��]���@ܱ�Woo+.�/.�`�mj������"�RA�H�dV��ӊ�!�n$�݂-�̍��غz;��:g�ɟHt���s�������WI�ͅ�tO��J�=�n�svq��n����� �yn N�����]���Z�iݽ8��7n��mN�z:��M�jb�ǎ��m�͎��.㳔��k;!�q�l�rz��k�N��J����wj�i�9�!����C�ݻ: �\'@������gc��ewdw7<��r�v��b��t݋֗�qt������bx�9���t�­ísA�n#��˷��?fY���ݕ���X�w���A��݋�ܔ��ũg<�7�1M�ݶ�m��t�Е�Y��Uy�ƭ��Kt�>뗪(m��v��d����+�V��@����7��j2��y�}�������8�z�������G6Z�"�հd��vd�[vt�t�玶�v�Y�i�oB$^j�[-E��\��Y'*6�y7 'kwv��,�z�� LTt2�yNk�,���cr��u��֨D��L�D��fK���oAB�x/����>j�7�[��-���;Nt�n�3�����1��;7WH�zL�N��y��±6+m�&�H�U+m���8�c�gn��ku��?#�Xx� �#i̙&2l�6��NBk+������tG�YCԚn��:�؅#�<Bf���ʏ�����-�X�1>��
�x$�,�C�� ��
s����=ƌj�(n���/z�d�ƀ F����9F�G��!Z�3d}��lm�Wev�R�1nGl�׬yQ���{�B��<�n�o,��;�&��߹ߩ��?^jH��zQ��g�ۭ��<(�ڋ@���I*CL��u���jё�@����lu|$(��Q���OSu,LDز	�y=
|4��Vh9�G��z�B�B��N{����m�4�«��	\�g0���м#VQ�
�����hqȑ�ޏ�x��<|����acNT
%lٿ��Aʘ��GݑV�N! ��%��ȋ?^�����cޓ���.ʟ��,Ʊu��O���Ђ��A�XKY;�/����y�UF����d-��c�I��P��x��ߺ�*K�,�V���� }�M�庮����O��(� t&3_�ʱ�!e���ۻL�Wek��"t�P>헏\�a������:�#��}_�?f�n�ʞ��&��!��sv�z� "\ة}��&4`�DK�� �bjG�I?#��M�$x(
��1h��͌�v��ŧ�<��_�q���r���9_rh=�P�e7<e� �{�CJ�M~ù#��B��"`�2����o��ĺj��v��L��1���J�����_۵�W;��'�ܠ�>9^-,�IK,N���6�P��/mnÝ�O ͇�3۬s�ކ;L���Q�Y����F��c�/RTۈr�f.,��H�2�;�ye#
��}q�մ��^|�h�)B�9DUiԢ��E��Q��|�}sI�ۉ��Fc0��<��q�y��9\�/���4��|���"}�^��4��\g�y��-g���lϹ+�j=�܇��I{垦��e!S�NBHQڣ�]Jf����T��x�K��b���7�B�����A䶆�ۉu���#���T��� �z9r'ػ�aL�
��<j��߇�e�n��/=D0R�_��T�����ڰ�� =���V8D)�Z���t�S��2��a$�P\�����K�`YUg.��ؽ����e���놤q���ze>Qj #����B��:�yk؄��;������2�Q�=�����K�R�y�����q��S��R��i��e��s_x!�	��)⇇%"4Gr�(a�]|ZK�kx����B8�4)J����j�fJg��}�I}���絀ǫ�\z>W���ǁ�9���6���È\��i*�Ԙ�QhqQ�g�g����+o]C�̸�?i�;L��$�lM�`[3�6�)Q����x��7�a�` �qX�}ՠ�5AM��Sf�I�'��������.��@���)hAO`�B=�����^�����r�3Ϲ���Zn��iQ����(��2G����G�ÒE���/�!n�L��ߥ��j�߷�X���mn��33Ɲ9�����d�Bu�����On�\��&E�\��N�>8݆U�c����������uʃp�v^٤�lζ7a%щ�}����"�P���-�H�	�p�|�M�Ê�k�QB�XOӽ���t�_��攝( |k7M_6}��8�më�_8����X~��ڍ�p ��H 8�_r�t� i�_Z�s�</l��'態���Nmm�ܖc�Y�{�D�2!U}�Y��jL}Ս83�,ډ�7��:��ؘ�,�1���CV���d*i��_�����Ý\�=�w�c�:2�2h|��73�}�!��r\�9Q��<'z��:�BS�}��i�."�0��=4��q?5�C>^�Q��p4��ӎ𚲢T:\�!2KW���)����+�������#��X�{�ܻ�/�#���+D)�H}��DG�w胐wf�]G-A�wj���X&<�jQZ!�Z*l�k����؅g�Ɍ�S�c�������=J>�Ea7�&Ok¢��]�S��T�n*��Y06..FhG����#�&�_z���t������y����D���t��l�-rgUDt�֔��I|qG*\�"�.Jj _����g�Kk�ܕ�/XN�_>:�5�N���/��wsؤ-b��v ��A�]�]�M^�⧛��Z\�I٣f:ܠ��f^ey��cY~�kD�i)ۤY̴���ëi]��#9��(�e��&�Sow�7.	�=�WP�X����	hܫܽ{��^2q�����mF�ȍ��"(h��-n8ʐ�ԭPwV�'�f��E��cmu�L�\��:��b����	��4Nᜮ��'�8��3��ԗnh&7���¼����Nj�ؔڥNM�(�A�)����6��#H�!�T��pj��[z�^Q���ǋ"��q#��r�=X���v�	�s�0j�WE�5�4,˰l���Y�n%�)�-4AlI�a�%'��_~[t���� )��W�Y�� ]ʑ�F��3��_,�Im�ݯ#Fd�kr�T��2ǂ����������c޽B��qIMv�Ǽ[�����u���*�����mM�8���#���o�ٳ��/��ey~#;oĖ���N,y���s���؋�~(��[\����Q��.�]�U���S2��á`���#xr����%ZT��`�F�A�TD�QG��
�� ��M��Z������1?r�<,�� C�}�a�3�!8<��Ҟ���iY3��+�g,*d2 >���a��	OZ�����`���$;}ܷ�BE�N���a�*j��?@� (�/n�h��Y�����*���mɻ^m��f˅��.����#�4�6�v����vࣝ�L�3]���N��_�~?w���^p�Q�K���O�pQ�pg<�i�U�[J��5�H�K(���=�:�6� �����)~���r��O����E�3#�+���^�jC��ki)��f�|��=g�=��F{��<a-��]�H��/�c���LXD;�e@NZ��2�������I8{�(�b#wZృ�۷�L})3;���u7�5rH0�/����M�D�c�ϧ�]r��~5�@n�|�sئV ���/L�<G����@"�����r
�dq��	��8g�>/6�@Ā%
�M��T �,D���4�ݠ? 4���	9��<&�|�����G��S؅�N�����N�7�T)�G�3��v*�E��l�1�˸��KxB��m7��W�X��T�;�|=�!P�&��B��o��b+D���3�u
�p��B��MFh
��ǥ�E���w�t���v'�B�����1��x2@��KB��S�����~<
r� q�]��!4j��z�p��Oч/;s�.���>�@�
3t	�~���+�dE&f��H���J^�k�t{�^أ���X�r&�pv��J��K���z-�镠�V��]��g9l��4�R�S�xg��H�W��x�=�"�"��� v��8��Y������s9�E��d��X}1�k�~�xlh�X�ؓ5)�_d�#��6�Q��[Z!��@�P��x�=����q��T*��f̛��c��5X�'OZ1mn
t;�����;d���wX�kYǆ���aއ÷���d��d�&�ũ�h��=�{9.S��6�������bE�0�G�����_T�� ��r��Ƙ��x]�b)��a�<3���a�h5�0:�}�ЅpT� 4����)���4 ,���X}��͋�Z��a$�(�YFp�d��5�s��*��u�׊�����|�u�̐�e�����B�ܙ
�P��ZneI�J��4���Bw�1�|'�
s�t�jge�^��q'�A�|gJ����M�-�#��|=o�ZE�=�ώ�̐�
�dxe`�5��9�
<�_r�}�Z���S� �OC���x�ݘmW܅uh�7�q4E�|&����׹���[fEDH��W��Ǘ�ciV�tWEf�>2�O����qݩ/�3� 3��ϼ|�u�Rno��xq�%�x�3�V��Il�jv'��Ht=�)鿕R�x���V8#<F�J����W�>���7�P%H��+� {�ZD�ì��|���kx�W������~���>���o���{)/�c�g�s�n����F��ߑ(#mJcb���*�:!Oػ����K�ߏ;����]�a�p�Ye%�ʋ)^�c�eJ����=~J�ᚨ���a*}}��#���[nǈ����r
��yj}�@{�fqH��
s������l{�=��_|�}��/h &5�ȶQ��
�!��)pN��2"2�BQH5ܢ�m���19���_K����43 �^��_]�ŀ:W�N9��|w�nJ�����<�hJazb�S.�m[����z���2�ܴ�9�u-����zw���.�W�8{��F6jy��~�YV��۸�zS:��o6o:|���Ս��ˇt��'��%ǒ�y�6{W2/"�7|�H��@�y�.�T�y�al>� ����?.T덭���n.L?�^�ڲ�j�U�*w�;��І�dg	;������v����|@�c��f���[��z닓�s?9�223�IU���d��4s�v؋��f��>jvv��v��J��ę$-٪��]�0td@RfC7������4s���i��[�'m�n��̓�v��<vN�ֹ66��S�Gu����5��۴Z;[��TJ��ɋmÝ��3>e+�N�=�C.�ۢ&���g�d���J�q�E�Ta�=qS�'+����P3��y�s��ӁwA��g����k��`����M���g��Fb^٭[����9wFt�ޫ�i:-rzV �M u%��g�(kz�wlcn;#�K��M÷n�{\�����>s� �� �]���y�<��u[�Ŷ�9��]gp6��/n5˨y�86�;��;av#��nF굫8�O�.���������Y.���K�l��ٛP[�Uݷǫ[u�c�r���M�8�y�/���*��]�~�;_ky>Pà噏7]�0���\��ǻ�y�ż��y���ʫ���Ƙt5�kX�Sz�
�J�T�xa�l��G1BH��fc�Z��V�݇`�z^�{&޻�6�s��ɡKkB��9:��������fN�Q��'}�GW�y�gFggv��v��Xg
I:�oZ�&Pы�v9��陲5&m>sc�%�\�����ϵ��]A67+��ܱ|�l��I=c.dwen���.�$B�}��.�9�ė>1�qq��ȷa�Vs�X��ǭ��n]�l�rv/X/;k��M=��Me��5~�} gM�
a]�� o#,
;f*����R��	2��\���B�{�}���4Þ��S�v�|�^�uZ2
��f ����r����Jlx�{�j9@ ��u_�e����[���+��;��$����/I����̵��3+�Cz�����-~4�����j83�ֱ�7��377����~�\�ᠱ��s9f�ɣҐ]����}Co�l�S�0eˊ]UJЂ���o+GB3\�~ q�[|+�����+�U� /i����"�����=�u�\�=�T,��NP�������:��U3��-�=����1�Pxb��/��?X������dm�./wټ�RY�zQ��"r/r4�$׿���C��P�Tf��
���}f�a*xq��R�+��F+�����m���8�R8]��4�&�(��H��
��s�)���h�y��.o�DDH�o����P � ��nl����8E
���x�->���p�VTOL��\s��{����˃������B���f���&X�7F����QJ�t���SZ؞�3C��� ��n����M�R�9Kq������Vq�~����ߐ���Ɠ_��
�?���"<=���О�2����S#|HS�=��T.�x��#��:e��a��>{�P�^��ե2�1.�~�o���?Q���r�Yw���z�6��H�m�Z��
�GL�bsb3u��yݔ.�����D�h��现��j� gS�k'�h�DD�Gm���T�t��٬�X��q��2�r�6�,�T앰����ʲ�����Y>�>}��ՈS}̀@Q���c��J��W�dy��5q�v��� =�+=
||=��`�|J��g�~ }�26�)�?�*K*;i�W$���i�Fm����We�/BR8����@��9�ɰ�#��J�1%8P_ �kX��i���@l��}����{29)��Ί��u�	o��\,3��6S���0�u=�I� @�J��Z���W�-9�������a����#��Q֌��Ս�a%,���;�_|(Ǽ7��C^(�Gע���YS��6 ��7�6&�E'�������}��2�fy�0G[8�ޟx���t����D�{��o�A5�=!�F�<�c�-�0ٜ�7�Zk��;�V�j��������=xb+JMy���(N(4�@Ţ'-���+�v�>�E;a��D�4���r����;���B�{�G--�y��a_��7��о�
�1��TFp�15�(��o�if�K��%�
9�0�M���T�3Y�.��]9�|�=������-}�pf9f�$iz�Β�j,D%m�����-�֕5��s��ƾ�~x��X�#5�ax��L]��/���h��&�G�f��8u��{O����u	����.��"Sư~�>CyoV�#���7�~�ENR�R�D�pm\��3��{喎q8�*�$М�<��+`zɮwE�u��W\s�����O/��'�ϧ���7m���Ry�]��s+�G;�ɀ(��!��}�?]��؛��H��z_�A�ZH2�6Z�ᕕW`���e�ʓ>���H�����we��3�����zVj���~����Nxx>[�A���[@�õM��q^#�}K��lC9YɁ���h����:��&��7@�d�,j�c�k	�dyC�E=�X�>�ד��+��ܡv#3�wIMK�3&�xEb|��ש��x��d��뀉WQ��R�@T�z�ĕ�%���|l�`����1�!����c�x_��?@�t�)��x}�Y���Ⱦ<(dA���� a�[�x����p��E+��B�'k���P��s2k���>�<km.�+�W�g� *�<Q�c��z����3|���k��tj2��P�7��c��9	4[���J��R��������e�W�� h�n�wE��ݮ�r����5���k��8���
p�Rgf9�v]o�sdj΅˧"��x��H
��y�f��~'wp�{|}�����oe��ڷg��5�4��j#X�l,���p�,E����*X#9On	gc�-�%u����J�[�S]+��2o05�sQWc��f0T�(��UV5D{E��R*�r��Ol=��JfN��n�w{��PB4w�:�mp�n�#~wR��_������W�J��a���=j��<�"�p��aӼ��?�e�y��g"�Lf�B�-���<�a��tc|\�Vn�c3�ӵ�Rt�"�Ml��r!e�����*�*��tW�b�3-�We�"���i�3wx��'��h���"��)�r��-7�E�#{�0=
�r��n�71oh��ƵPV�H+�;� ��z�K�ˣ�l������FX�N�sBX�;n�Nj���
96�^d�����ܯ�t2WE�9o^�N
Os�Û��κw]sx-��m�h�D�Uۘa6�6�����\�<��wMA����?���0z��^E/�����"��u�?�q�����q�����|�O�KZ�X�,�ʨ�j ߼�ė��g-� N�T���[�<�G7��xRa�܅g�9n���$g��}��B�G��.�~u�c+=qv�m�����a�VQ?lt�^+�캦'��o%�[Qcf|
=���Y��&�O�C�i||�Y�߾B�<�c%%N��rGY#,Z�31jGb(v�!ᰫ�Vg��@��<�c.�yo�m��)�0�%��9=���7�@jr���T�C����ߗ���"�|gmD���hf�P����ܚpdٹ6�,;I,��。2�B��秞��3N��t!�e6�Wmt7S�m�;��`ֳ�s=����l����9���=v-=2��v�o	Cˊ�=ä\��9��΋5/�Q��n�3���ȇh��Ȥh�����`L���0��?x}��V޼����c�zn����j��7��g�!��N���js���5v�@/ �E��BD�<G�Mf��{����emU
2�LAe��x�L��q����>��GGkV�s��<���h��Įc��]a�9�ܝ�1��e!�X<�.~0����յ3�l�F	<'VB��{��Csܨ���'��e�3~�w�Q朏/���C�D_�x��a��7���w�����������-��Y4��5U��55�G� M!�\� ���\�>s�k�}�뾿fɧ<|/)���F�O�!��p�ߢ��Y`�&�"t����"&!����`�^��� �3�[�04�rpx�)�pW�Zߐ�@D��1�i����f���jZ����>�����Py
{�>-a�[���,� ���j>��ܬ�=,է��	S���1<��R3���D�����b�E}���!Q��w��{0G��{O_v����
)�[��=�{j���(ͺC�uno,���� !ᖠ�z�n�u���jI-N�v���3Y2HS��m⿦ 9�^������'�x	���F)����S�J����)-̀@r������i�첓&~�4I����F�+o�mǠW�c�����U��Aa7{�֝�T}t�fq���?Y������n2��]�5���5��s9v�,�<��n:>�q/��W���F�[��,��1�7����m,�?0����!E�O"�7+-f�ٗm��6�b�5T��%"!�#�L"���*/��q���Pv�~��@�V}�H��7{I��qL��5����wKp�x�6\�3C�M'�8fqXx��O�3���9��
�N!�FIPWI�,5��2��t��� 1"~�u���d���s
{��JdVi��Hδ���*�;��*vX�B��2$JI;�(���� (���?	5 V���3�,9&=зU}Λ[�&�^�XW)�����N�J���m�$l�n��*��.X��V&�m�IZn��2k2����Ύ?	.ŏ�v�[d�#��ޛo�������)��lܮ��s�s<9�����I҉�ۘ����9<�����#SH�:�R*��{�\h���h�S~��<0��=�`�i}:��\��}�=dG,��e)�A�
�PV�o9��&Er_h⏽�|�z��䑙��F9=�����l_���R����&� ��U!�+�lI�;���^| �O��r[-L�;,���nd�wn�
T`&ɾ�y�$W���E��.J@/��f��ӆda>>�mA����＾�F�B�F�vڣj`l,��fH�Q+��c��]=��=��Ru$ �=��D]}��`#�֏Ǩ�~�/G��ʼ@�\z�[������o7K�|���o�����>�����UT~�8f��������Ϲ�o�?&:�t��GG��93r�q��^:\�/���9fٛ��u�f3�����M������s����3���<fΫ��]g-���$l�g�m�&� u�lw��c8�����6fٕ�6�gN8yx7e���<�g0�����sӝ�=����͍F�
ٛ6�ң׎��㗻���?�����{�=_���d��3��N=����l>��Y�ۣ�O��韇�����{=���������~w���}�����=�}�>�c���}^��vy}�{�l�9�}�>���������t���1�����[a�/�J�����~��|<6�Gp����M�=���7��w��}�{�����}�����0͟��o���������k=�_���I��:Y����4|��7������6�pz�z���÷n��5����_:w�}'�~ߑ����s����l����Ӟ�����<��$B&��d[Ye�&�,����H��&��E�Z,��Ed��Ȳ�E��YdZȊ,��Ee�M"",�k$k,Z-��"֬Yb�i���"X����bE�YYY"E�D��%�+(�VՊ�j%�++H����Qi�VH��f��(��H�%�QX��K+$$VI������S%�+$+(����b�Ք��"�1BYY��-id�Q,��F�ie�B��P�VV�6�jąb�+m��Sm[`�6?�6q���aLՌ�5����f���E6�e0�Ք�H�F�YF��X��AYYMY��V+(���Y�&)�K(��&ڊ�[(������-b�,Z+$H�j)�����YBYh�V%�V)�
(��H����Y���(��X��,�VQ,Z�"֖H�VQYE��-Q,�ZkY,������Z�"�Y���-e����"Y-cE�Q[-f���V-)��YE�-Z$KkEd�e�ȑD��,�[E��LȖ�\8kE�Y2k$Ye��h��Yd"�Z�"�Fȶ�,�Z-��,�dDC,���-"�"�&���k-Y4KE�"",�`�h��&�,��k&��Y���B-e�-�l�Ȳ�D��D�DX�h��[L�ȅ�D�Y�k&��mddF�d[h��h�&��,�m�X�"���bȋ�,ȶ���E��l�&����&�Yh��D�,����i����2-��Ymd�b,�-��Dh�Ym�5�Dk&Z�F�"�h�b-�MŐZ"5�"5�"k&�X�,�[ZœE��Y2�i��b-�L��-�l�4M��D,�[-5�h�d�i��E�-�b,E�2hE�&Yf�md�,E���["b��ɲ-�[Y6��[-��X�["�&�,����YlE�XY6�5�"��-�&"#E�ɲ-�l��,"Y��Yf�2�h�YdL�D�#Ym��X�m�4F��M��dȶ&�h�dh�Y��,�LDe�h�E����pga�l��k,����FE��M2-�-���&�B!Ad�Yf�,��fYm�mm2-�ml��h��b�&�"�d��,"e�h�k-�[Zh�dțYl�dF��[Y,Z5�Dh�,E�ɴM["�l��F�e�2-�Y��5���4Y,�E��h�L�md"h�e��,�DE�!kD�["d�E�bɢŒ��l��Y2!e�-�k"!kk!��ȱdE�MȶDȋ,�X�"MhY�e�Z�Y4[D"�,�E�E�Yd�h�ɖ�,��Ye�h��Ee��%�E�֋DMmfyuv��M�'��qr�w+�v=�s��ǧC�6�=�6���~����v��=��?�g'��?ǣ���q췭�n�!�n�s�c{�7��������߻���/���w�نl�w�g��>G��=~������������{�?������}�o��_�]S��d�ۧ��$�;���������?b��a�>�ӻ��~�\���/������x��^?��~��>sOˇ���/=�f�l�p�F�����e��_��w���g��ս��q�:��O����]�����M�n��U�.~?���:��c6[#G���~'M�^̇�K�[���&�]����{tYۮ�;nx�q::7c�;�pwo�wf�������>O��ؿ{��^_�a�?������,�w��w����yg��}�w��m�������>��3�������|���n��b����Z3���]ñ�ϣ����:��f˟���S~��_����0͜���\?�}g���_���z�v?����q�ni�}3����7Lp_/��/�;��}g����/G�E��=[�{~�>��;v�i�xs�������/_���{>~�{�����^p����G��l�g��tE�~�����������z��}�r����ۏ���4{�)��ݾ׀�����9�����?k��?��)��;v-��w6�l����-�gS���:?뻌����߇c�����z>�l�u�p�DO�{?�.�p� ��|f