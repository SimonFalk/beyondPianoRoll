BZh91AY&SY�p����_�ryc����߰����a�~BU�                          f                         !                          �         �                 @     JQ*	  )UR(64�@4Ҁ                                                                                                                                                                                                                                                 Y BT                 @ 
 P
��4b�` `M0F	��� 0�2h�14�@��`�M4 a2dшbi���4�&&�h �MRIO*{Tͨ��z!�  2 �
RBL���	��J~��ji�OSjlԛ�U0AMJU5<(z�  �M4C�u�z^��{�'��i��O"*���=��
���`�RܩQR�T�V������-�1��U)NH�m�L?3�?����m����i;XFYa�\V�Q�e�m3�3�ڪ����a���U)�2�`ʺd9�12��rN�V�(�aS�T��^��<��6?��������ϗ᾽WJU�¢Y�I�))��)��f�X͕�̣6S[:>�=~��u߱xf�yϹ���n��R������cG��j˱�����u����xc��Y7������m׶��=;͖�������nc�V�]�\����B�J�X���[�l���jS�\S�m�������p��n5�0����-iqI�%JC����Ꭽ�)Fζ�P�b�Z�����y/%-��$�Z�ڞq��1�8�5�Z�T���:��qıե(!I)Ŭ���18��Y�:Ք�Î��-LZV�imHk���:�B��ia-�p�-�]K�q�֗J�����hcY��:�1HbR�t���8����!j-	S��C�m.6�1%�,b]mG]pRHqDǭ�)�����!iSjc�c�!6�m��l%�����b�Z��kuũY�I�qjB�KoC�V��<��B��]u�1�RP�m*SqS�z��t��K�J���[�:ġ�6��*C�JP�yšH6����ڞB�8��!M���!�hu�1hm���=���:���(tm�[ͱg�����l[�:��uLqhqq�RN-im԰�6�]!*S��=�1n��!KyLb��%'V���Z�m��iK��M�Zǵ�-�1hSlJ���m(CjB���!M�����qM��Yhb!�0��uN6qŸ�یuN6c�{jo[u�Co!m��yib��!��un%6���n �6�kJ�BR��n!t�X�6�5��p��ĥ�6��Cm��X��a�����c�����!m�����ڒ�[�ۈm�cn8㎬�����:�یqL[�y-�m1(Z�-M��B��kmM�hqG[m(mm����š-��IŽ���<�Ju�Qe�d:���!iQոŐ�6�n:�C�--��[BT��n1���Ҷ!ip�I	K�3^q��K���:ٍ��Lq)6����%�q1qz�Ԅ������c��J��u%��1��֤�Ÿ��YkKo%��-�,m�%���8�[C�BKqIj�yHQļ��uJ)iS�[[qmq�c�mM�[jZ�c{�m�y�]ym��Ե8��-+cΩ��6�ĸ�-+C�m����l���-�	m��jbX��� �R���(�N��LB�R���K��
m�q��K�)�AHck[����mq����S���u��-K�,��uı
6�Z�8�\a����AŶ�J�8���T�)��m.).��8�!iF������ukmN)�m�:�8��]R���+BX����m+J��%+c�R������㍺�X��Ԕ:��kR҅�IJa�%�6Ķێ�uM������ťu&:�Z�k�[��+Qe���ĥ]u�Ѕ!�Ki8�u!�)+B]m.%iq.��:A�:��ZXZ�qLq�%��]um���q�j�q�lA�Җ/m��S�8�ַ\Sn�it�Ї\ZK�m��1�u����u��\:�P���!H�]RR����mm��S�RP��-����XR��RV�[f֔1�-�t�PJ�Yn��Z�J\R[!�[��N�n���l��[�))Z�:�X��ciC��K���%hq�)ic����R[Z��!.$�k-�:�hm�8�ͼ����6�:��qKi[B�R�YN��kq�%-�\q�-,S�m���C�c����JS�S����.!�b�uIa�%(Bm�%�R�ZX��K�Y)qLlٱ�t�uM����P�Rպ���8�����S�c��M�a�l�ҕ��8q�8�ciqN�.8�c�q�BVm�m�T��)n��q��-�J][jR��[q��ږ���1	:�1�c��R��R�-)�J�A)K�ե.��:��[��uZ�S���[u��R[q����m�8�!���P���i%�R�!n�R��JRS���Xu�:��m)6m��ť�!խM��-iq'���!�mN���C��ĸ��6��u(R�S�S�u�H[�-�q�:�-�!�:�6�R��Q��ڎ�[qi)(m�1*K�SJZN��B�b�p��ۄ�R��)Z[u
u��%m.6�҆��mlJ�J�!�V�����n��!�6�������S5jRR�Jq�8ڔ㮭lq�5�-M�R\8�
6�\K[iBT�-��l��u��uթ���1�u-���8�1iSfmÈm՝bַ\K�b�ű���jA,K[m�8���)-��R��i��	aIq.���J�ۤ��A���n%�����aĺ�%N�C��u�%Lqպ��qԸ��Ї�GQ�l��[�Z��ě-,u�A��m�;�ۯ)��6Œ��ڛ[n%M�Hb�y
b�B�ǥ�8㎬��%ǝa���--��X�5D1�-�Ӯ��ź�-��ӌB�m�!-����Rؗ]q����J���uŰ�T�B��un��X��6I:�ke�J���Jy�!屴��R�C�q����(c����m�-bV�R�����|��-ҜZM��-i���--�HCًm(:�e!
yź���jZ�mC��S�mR^[lu
q�%o),u�%K�8��bZK�RV�]m�LJ[Cm����B֓Ԧ�m�.��<�1.�Z�R��m��kic�S����Ŷ���1M���K���-d�����[��ěq���[k).-ĥ�\Bз\-����[��ێ��lA'N!�6��Ӯ���5�X�뮡�:���,�SAjq*B�y�J\K�Cjq�-�!I8���[$�1(q!��^կ]C�Z�Y�Kǒ��)�<�1ǡ��ג�m��SkC�1-m��6�	bT���1��[��H$���yz�-�!ӬK�)hm��Rإ!.!N��ض)�k��αE�G�cC�:�V�6�:C�u/u�:K�q,<�����8�iuk6��Iձ�8�1�:ۮ�e8�iclmn8�hb��$뭱	R��\Z�Q�u�8�o%.��Ҷ%�y.%������q�\�oi�ťèylR��IIS�-�ڐ�!N;N����]C�Cn%y�Z�6��!��u�!�ĩ�:㭡�R��JHK�c�C��ٴ1Ķ���4�BPyd��!K�b��RB[F��B\[�1�՜u-��V�T��K�c����(�:�%��iqlc�ZC�:�B��bئ�����mJq�R
m%�HCiqn:���M�����ZChu��J�c�S�q�Ц8ZRb�m�[b�p��\uiB�q(b�u�%�6�!n1���Җ%�ی%�B��<�XuF�l�[q�:ũ�-����kq�8��m:JV��{�!�yO1�<�)�$�qG�(�6��q!�PǭHZm
u���^CV�X[X�!�B�ۈS�����8���1�ҥ6�)n6���(�mԱ�j��%ǖ��ġ�C�Jͩ%�!���-��3V��X�j[�A��ىqn��8ۋB��+TuN%�KlBV�lm,J��[6ԥ漖ִ)��{�����%*!N��1.��l(�mhmb�҄%m�m��bۮ!�uJChb�B��m����Q*um�/!o<�J�8qN�qj6�8�hbͶ��&Ԕ���m�����6�Ŷ�+u���)պ����Ԗ%mS�V��K�[���Skq�%�1��[�mպ�5km�p�Z�RV�=��:��Q(B�q�Kn�kq�!.:�R�c�c�)�J�c�������R�8�����).%I'�d<����q��X�Ԧ�؄:��X�m�����mIc�R�J�[K��N,�!նR�㺄=�:��� ũy�����l�X�(�-�q�m�B�� �\SV��Z]mR��VRm�%lkC1���]m�R�%�!n-�qu.�8��K�cmhmí�ĩ,uhCm��JV�m����1ź�X���T�<�T�m��Ϥu��.ks�����'99�<�s�R����k�����f��x�L��|�ލ�m�K�l������Luk��x[\�^�Ե�8���)�d��[���������ם��]�c3��;��e����2�r�2�e��"n�����W*�s�������)��AեK-HJ�����T��-i!jP��kJI%H-IAIBڄ!$�HB֕�BT�-*Bҕ��	%IJH���ST����)Z�B��!	BE�%E-*Z֤�
j��)KB�JV�(����KJT�))Z�J��%-�-HR҄�IIKZ����%IBR��J[P�R���J��%hBT���-(Z��ֵ��������R��Bօ��RХ��R�)(B�!jR��%���
AKQd��-hZ֥��c��J	R�PBZ��kZ�)KB�5(B�PR�5jJ��)IB��E!Ij��kR��Ҵ����-D�!-a)R�%JJ��5(BR��-IQD�(AKJ��!HJKRJP�(���������V��B��%HZH)JR��k)iJ�JR����iBҥ�HZ�--ZK!k �)e�KJT�)+B��MQK,�KAj)J�-*R�j�K�-jB҅%CP�$��%-ZԖ��!KZP�T�%)@�-Z�B�Z
B�+X�-*R
J�ZԄ�IQ*B���%%)J��-j%D�
ZJZ�!KR����-(Zi+R
BԔ-R��HZI(��*CP��h$�����)JbR�)IJB��-(RԄ��!R�ZVZ���)!hY(YkQKRR��)R���KJ��)HZP���%$)Rд�$�RV�-jBJ��JZ�%IBBHJ�Q)Z��JЄ!e-IQiZZ�b�-�B�Ւ�����KJ�!JQISR��	QiJZP��%HB��)(ZP��+B�R�)hR���-(B�)R��Ԃ���BP�%	R�RBԄ!KR�!k%	B��V��Ԓ��RҴ!mQRP�VJ��kQJB�)
Z�-)Z��T��-+I*J҄�Zֵ��%+JKRHQKZԡHRV��	%
Zխ���)A)Y	jZP��KQjR���KR!hR�KP�!iSV�!d��%E�-K)
[V� �Q
JT��J��KJ	B�!jZHJԄ�kRR��(ZP�(��%(B
Bԁe�
!%�kZԅ�e�
QJ��)jR���lb�����HZP��d�HAIBХ!SP�-jZ�)d�%�jBT�)*J�����
YZ��%)R���R�QKZ�,Z�����)!d�)YKBR��Z�Ae�HKRRД������KR��ԅ�jA(j�RT��KR�RI-E�Ё
J����%+R���JZ�-)B��Z��!ZV�%)ZJ-iKVKR�!
!iZ�RB
Z���YRRR��iQCP��$�+B�JTZV�-%�iJT���HKV��ZR�J�%D�HR��)JB�CR�)+J
Z���jB�ZHjKJV���	-�!)Z֕ �V�-IJHBZ����-IJJB�!jB��)JB�%Ij�!hRԅ%%-	R���mZ�R���hJԔ�kYJRRҖR��%+R��KI-(RY5
Zԅ�HB�)mBT���-)RP��-!iZKR�I�(YJI*J�եiR����D%hBP����)J����,��R��kBԵ,�!*-IZ��,���IJ���%J!iJ�R��)E!BH!(J���!MR���	)(B�!JJ��)!
)KI	RVRҢҴ%IIe!�SV����%)Z�� ��
RHjV�)*J��Ե+Jд�KJ�҄%j-K)$�(��hAd%*-B�JVZ��*Z��$��AkBP��Jj��%(-kJ��hR�-K$��E!*J�J���h%�-KBւBT���R��%H-hj�J�)iR��%	JҴ%(BR�%iBKYk-%D�e��%kR���jZ���!MAH)hR�!e�jSR����)MJ��-	Z�,�-B�YIZԄ!kQIR��!IQ
-*Jҥ��)iR�����K-jI+Z��jJօ�-BҒԕ�jRJB�(�%+�-J����kj�,�-
B�B�BV�)d�Jք�kB���B
I+ZP��*RB�QhZ�!)B��(�����J���IQ*Qh��JP���JV�!jIiR�R��Y%��,��)R�0�,�T�)
Z��)	I+R��JB���+B����)	B	ZVթ	B��%JR�ԭ
Z�J�!(Y)ZP�)	ZЅ-+B�B�%(B-JRҕ��(�HSR�!KB���(��	Jք�iJ���!kQ��j%)-kAd�-	ZV��)AE�iQ*Z�-	B���
Z�Y%�%(��(Z��
Z���J���J���J� �-jZK,��SR�)%!%�+Ae-�BZ����BHJYJ-JZЄ)IZ�J�ID���%hJVR��	R�AKjR�-)B��Ң	)+jR�-
ZJP�$�)Ij�I[Z�%��B����-d�+K��k%D�d�iZR�!ZJI+RҤ)kJ���+%K-	JЅ�B҅%kR(��k%R�Bԩ
R��
Z���IR��KZT�����ZP�����Iij	%K)IZ����R��� ���Դ�HjV��	ZԴ�YD��YBKA(B�!iBִ�	-����-+Y)JТ���+ZB�����IBЅ���-$�BT��)I)HR������Z�!
Z��P��e-JЄ!HJ�!%%D����JJV�%JR��)"�RҤ�J�ZB����)hR������jAe�HR֔��-ZT������BJY(BV�-HZTB��!*Z�%(B�Z��%kJ��J�-hJP�T����Zֲ�����	BЕZ��H-kB��	YkBTR�)BX�-,%
B	I�JԄ$��KRT���Z�B�RAH%d�I%iR����Jҥ(��BR��	R����Zִ�IR����B���-*[T������,�1)KX��$J�!�Z�)*Z֡IR�Z����K!�R��D)HRִ-�$����HR�R��iBԤ-E!YkJ�� �,�!JJI)B���hB�BTBԔ�Rւ�)	(�-KB�J�IHZ��)*IkBJ��%+Z��������%*R�)jJKI
BҔ%KB�JT�(����%�h[V����KRZJJP�-E��iR�Z�B��,�T��hQ	H��mI(-)-hb��l%(JP�)(Z��kJT��Z��kQIBTRڄ�KZT��*Y$��)kR҂���*BҤ-e��J�������ZB��-hA)B�ZV�T��e-k)HCP�%D)+B��Z(���KJ%+%KZ��Zԅ))$��IB����-kBP-kZ�ZR�)�B�ڄ�������!B��,��hƛ���5図n9jm�m��po~�%Ja�\�z��R�鮚箍�g��q;o��R�7��̱���T��Q�?�!������>F=����?Զ��BJqť万X��C�)!���:�n��m,1�!ҝK�ukB��y�J�c�y�[y*qy*y�mO0�q��[�1�T�1n1�Kn��6�bPbV�<ۄ6����:��b���!�-�<�V�-ג��h:�ka��m��0u�Lu�n:�:���:��␆1*KǛq�C͡.-�:�^)�T㮱�!�%�ꐷۋb�So%�<�!��Kq(q���T�h[kI�Sͺ�^BXٌx�[�K�%��K�)OKlRu(qCۮ��jj)�6��q���BRǒ�)�u-��:�Z���y*q�8[�[�u�:��y
K�Sm��\[�ygR��S�co��Siy�K��S����Z��<�֣�miR��V���-���kb�J]In����n��N��JR�y(yg�qhp�]yť*c��ǎ��Z1�6㍼��mn��ζź�㮼���LZ��[�Z���%ĥkm�,�Kf�㍼p�K$�f��k<�R��S�C�S��+0���n8t�o(���ug��qN1lu��6�1N-K[�K�I�0�bbp��R]R�[��An��6�b�c�B�BV��q(J�Ǎ�ǌQN�Ժǝl�����[�Z��-ŭ����HR�y�����,��l8b�!�y���CjBT�).�jC�u%-�8S������P���u�1�-M��Pǜ8��mKQ���
uN-)�<��B]RG�y�c�)�0�8���խN$㭺�R��Kn���BK�:Q��-��gM������]c�B�[S�:�ͼ�<ٷT�^:����1�)�KhCn8�8���q�b�yIC�<�8ۉJ��!�y-���[<�Tű���u�C�hqIy���!JR��yԥ�%�ui6������ոڐㅺ������S�SΛJ���ۮ�����m����[�CVǔk�1�Ҥ��KlC�AiBC�u	Bu�8��B�ռ�m�^q�uk[�JN���K�g��QN!�y���$�҄��yht��8��t��g�qIy��m��RJ)Ky�%�qn�c��t��뭞[�%�Cά�:����.���KRuE����6�SkR�q(u�PRP�<�1���B�C����b�뭡B�u(Zև]B�m�ŭ�ju�-oCκ�����؇�C������-��RXB�%n����yԼ��K��m:��S�qo)1<�n��J�ǝu�)ku��ΡM��6�!,c���:��1o1�~SyM�(b�CK���S�R�p��۬mn�⒇]q�)��[qlJ��S�Z�m�8�S[�A�m�KjAĥ)/-�[m��������R�ZN�ێ��m1���J�Kn11+c�:�1���c�8��!,j���1�<Ǜ[�6[c�u��:��<�%��hp��<���Vm-��mo:��u. �6��-ձ�Sn)����q�6�Bu�y�8�o[kcͶ�6���Q(R�bq�8u
J�Rα�N%Iq!�u�1�y�n��-�u�μ���8�1
C�u�SkY�m�q��ż��ۈY�[S�u�-���m�iyIy,J]u�8���ֳ�A���q�)�ky/)op�-M��8�o<�u�P�%�<�%*q��<�-O:�P���� ۉy1��m�)�^uc�kb�)ŭ�m(mo!�:ŭm�,S�IjKkJX���o6�I%mkm�yN%���Lu��S����V�q�1	RX�8��CkyLKiu�%�y��B<�\[�R���8�$��)�Q.��[�q'�S�m	q�6��K�u�1O8�-�b�8m�P��(t�u������ה�ku�^mjSg���:������)�6Z��[S6�!�J�%����!ǞC8ێ�*R��؆��^b��J[x���:ġ/�1By,b��:�Ԕ8ۦ%�����8���RS[im�J�q�)�l��JЖ�u�P������1m�)qiRHC�1Ip�X��Bԕ��%�<��u
m���8�%�	y.���m�8��:׉yĩԺ��b��c�c�:�!��<�q�:㍶��Rq�-� ���1ǔ�8a���1*Kj<����6����ZR�R��R����:Q�%n)LZ�uĺ�	y�ا^Z �ͼ�%n�պ�:���R�R�m-���%ě[m��q��1G^Byn�Jan���Sn�Cjm���y���[jm��q�^u���m��Q�[uĭcn:�%jq�^C�)(y�y.<�u�������p�:Ķ�m�+K�mF�u�%�%HS�q�\J\b���C�-N1�^uN%א�c������j�K�8��K�u�����Ck:����.-.6�u󎠧��mJ[�y&6�ZR�[bm��m�X�!RR��0ۮ0ǝmN1�HmJRێ(��[��-uն�x�1.���u�!!�R]b�JIJ[Ω[�q�:�\y�1��m��qq.%mIq԰���m)ն��ڞy��[K�Z�ml)�	S�1��҄���m�A�^Z��!թ�����`뎩.:�����M���y'����%'yטٴ��V���]c�ձ�ĩIy�J����T��u�u�.q�K�yku����P�F�C�K�ckqy�!�8��S�)n%JK�[u�:�RV�yԸ��Z��l��[����ǜm��u�[a1n���a�Ƽ��q�8�����%Iu)Rcn�)bSf:m�t��).��:�S�S�!���c���n�	qġ�0ژ�).�%�hqg�J]m��!�6��m�!�,�P�n��S�8m�)��chC�Yא�-�mԥŜSd���/!�]mSkZ�m�Pm�bR�X�6q�)�mեպ�ĵN8�[u���ĺ���<��T��!����CK�lq.)/)kqE<�!lR^%O:����1�cV�奵�y�Νu�C\8q�o6�S�q���ͩ�[
C��ǘ��uM�luM�S�m�u�S��䶖8K�%D�ǜ!ǘ�Ckb�mũԭ�)�)�6�8����B[u��<�^u�y�5�<K�<[[b�Z���n%�yԶ����ZZ�Z�SkS�[S���-yq(y�ź델�u�K�8�(�:��6��)�-�qǖŝq�%�k-�N:��:�hK�iy�K��PǜS�8���-:�ҥ!�JZ�[�q�-�-��8�SlS�Ku� Ŷ��A��qcK�[m�:���-��ͥխ�[m�-�<�ͩ�-�yu-���yn��ش�l�[lmgC�m*m��-Mm��A)!�aF!�]S��Ė�S�m��lj������n��Cj[�C�u�����n���y�C8��)m+c�)-��R�d%�N:�P����8S�qN!�<��C�m�N����][m��[J�Ķ�B[km�<��%�)*qKmמu��-�ԓ���έ�6�%��u��y���R�%�[�qO%����-���y�<��uIZT�R�mJ1��-�Co6ǎ�/-l!iq�y�V�u嶄��^a��B\6�kZ�b���x���j[�Kq�l�\m,uhm+Sq.:�C�6�^B��mռ�ַ�1�-�<J���Y�CkS�<���Vĥ��<�,���ڔ�����!6�)�^q�Z��.�RJ����ŭ/:��mLmԥ/~� �6cf��k�+�}�|Y>�j�'�ϟa��e��Ѥ�����=���s^�qb��ֱޫ���o�!��oQ�2?�P���z�k��b�BP�Ф��)JR
Z��Jւ������kZ�)jZZ�!JJ�P��R�J���MYj,�%*q�B�1ZKjԕ�k)
BЂ�� �)jR�ZT�!	YHYe�[R���!+BҴ-JI*!	B��!KJHAIj������+B
BԔ�jjB�-*JV�JV��+AhR���Z��)MZҔ�Zԕ�����!iA)JԢЅ��JR֤-JZK-*IKB���I%hZ�Ք�5(RPAk))B҅�Bԥ�hAZ���CV��iR֕�d�����-JJ�R��)Y*(�T��)jZ֦���!hZ��j[V��jJZ�RPRҤ�D���-jI
[T��	Y	ZR��jB���JR��R�-iB��!(YjB�!�-H)(Z֕)KB����� ��IZ�J�%	j҅-(JP���(R�(��(Z���(JRV�P�е���%�(Z���HA)!
R
ZP�!
J��HJд�))$��H$�%)J���*%j��II(B�5EJ���ZRը��*Rе!)J�%$!*ZԤ���-$R�JP�5$�)Z�B�A*j�ZJRҤ!)j��)D�E-h)jJ�AjZԅ)	Jִ!k-(j��-	B��-HR��Т҅-J��I	B��k)J��QR�R�ZҤ��U�t�.�y��[��8�o�chK�mm��)���%m��]JԵ����6��K��6���a��8S�:�<��VB�by
J��ԇ[%(m�b����B�uIy�!�ǖ~K�[hq�<�<��ѷq�-&ߒ����)��V�h~c�\S����^mԱ�\q�<��N��!��b�y�6R��\q�8J۫<�1-�R�mJX���}�m���-q���uhK��-)[��C�j�l����m����m�-1��qJKo�α,a�1��H!�Z��)B�u(q��������,ĸ�]mM��<ڔ�ζ�1�b���q�%מc���%JS�]u��y(m�-�Ԗ-/%.%��)��Q/6�J4э9��n8���%IBJBYJB���R�I
J����hJ��)-(J������J��%HIE��KBR�J�%KBIjV�--(J�R�Z��h-I!-�ZR��kRԄ���KBҤ�*I�J�!IBZ�Q	B�����⒤��ĩ��Y!N%���
uISP� ����!j�������B��?鵓�sx0���ݎ�V��?��]p��/���m'�R4�j���\S�(K��6���֦���t��������ڦ��P�?1��ZR�%�m�k�$u���'������cPy��B��,�Z�%+RJIJ�B���T�P�ԛAO��������)*!��%��c�m([�:����-弗^<K��b^[�qkZ����R^~Y����(RSlcJ�R���)�lJ��P����m�qIK�(�C��)�$�!�������6���	3N���8�_�cZ�n�G�����?8�5��~BPY��Ρ������MJV��)HRҤ�%%+l)lZT���R���k�I���Jִ���J�O?)�� F�o!��:�-l~{RťO�)lb�~u-�,m�lKg)�H~qg�m��P��	%�-����!�eX�:q&AjKik���1�-űF)�BT�!JJ�ӯ�)
B��Rд?? ��丆��cV�(I�0���J��8����4�
C��X" ��\SJV�!hJZT��$)	R҅�	ZJ���
JV�-kk�j�Bߘ��RS�J_�B��BMCM������Aym�hB҇���$V�)E!��P��-
c���ީ���u��y.0�O8�<�V���:ż�:��s����<��D �%m����Ҧ�Z���	m%)mMSKZR�8�^A�~B%+:��9�Z��u���j_���	B���kB���Ԭ����%��Kbҵ%~F�Ŀ?%��(jybġ.��6��C[A�C�iu�$?-��8�$��~I�HA�iHuԭiy�	t��j��[B��ƠqԜ?6~%�0��i? �����K�Qn���S����<������1�y�
[o:���m�/�<���hyǔ��8�\m��ZR��	J��+Z�)e�jSV�$�-(B�J�R�-d-!)R����-	RJڢ��kY
Zԕ-ij��!'�T���BRR��������
-	%iZ�JPJԕ!IQ�JVJҕ!IYIJ�YjZ���B�Ry�)�a	I�!���)�Y��8�X��	B���JRЕ�kB�R��,�!Ljе�iBҷ�%����SKI/ϛq�)+R�C�i1�~B�K����)�-k? �6�	i��AO�Bߐ�T�8�R��,[���bu���+R���]i���bR�m|KO%��S������iBJR�B��!KZ��8�i,ZX�-~u'K�m��Q��ĥ*yA�:�)�q��b�m�-H~qf1�%�<ű����0�Î������B��%M��:�-#h%)R��qmK�JP�X�)8ա�ĭ�/ǔ�Tӭ�%ǉa�1�q�j��AN%�B��R��.6���I��RMP�?8�-����? �������-���~R]R���+R�)kjT�вR����-(ZR��	C�󦩽C�<�έ+Q,~y�hE����mHR�����JC��LC�8�X�JClco?:��:�m�8���N��C�y�ߜ[�u�j�6�!&Ե%��l� ��ZuJS�ice81Ժ��jRT�R��]KTן�~A([Z���ĥ�]!H1�.����q�J��-Ԕ??x�RBRIJB��-%�RZT��%6���bqığ��bO?!%n��[B%�m�����O�ζ򒥔��-N��X�J��~6�ҥ��Rk�C��jB�K�o�6��Kyb�C��J�~S�JP���޼����hIJZ�(�(󍶃�T�
mhyM�,B���m�K	b^ShBT��\S�R����c����mr��kJ���J���HZP��Z����jB�J��(R�Z��������y��K�-�?%��5&!.�� y��%N�h<�\m	CZ��%�Rq�m��Lu�u&k�I�yu4ڒ~m��աIV�6�[ �!,J������͒ێ6��u�c�uJm����8���J5q��[�Q*S\�_-
u	R��5�e��ZRZP�)*Z�KT�ԅ-D�iZ����!IJ�Zօ�%*)JZ֕)�RТ���kR�j�AkjT�%h-AiJZ�!
!iZZ�5	[�I-+K���%iZTCT��kR�)j)HAKJP�%i)J?$�6�Ԡ�(�!
Z1���K��X���1e�Nb�ԝY.:��
J�Jҵ��-
Z��%	B�y	Y+bЍB�y֗_Ρ�c�f����%�����J�~K��P�ږ��_�Z����R�����B_���JqR��͠���z����[!*qim��k�8��]K��kKhG�:�]JP��B��ZԴ�jB�!D�
%+RVJФy,B_��uԜy�����Bp�?:���%�T��!��K�%mԡ*~~[[��o-��y�:�)���8��Jض��K�Y��HA��Km)ZqD%䔂\y�4�k��N)
[o�m��m$��1���R�����
b^CB�I���)�-hY�u�%�<���0�.Q~x�-ij�J��-	IkZTJV��	R֖�S�1jZ����������-(C�ŭfߟ���H�	S�ZԵO!�qٳ�ë�G7֚��Y���z�vc��?6����Km���n���Jc�-�-Ӯ���/<񴭴1�^�Y��<���8�Μu�뎡�[ZcK�8����yn��6�8Rߒ�͸��m�1���y�6���ly�ĺ�0��Х:�0���n:����[�Z�uKtŭlC�%d!�)O)hq�1+m��)uז�μ�-iq�Rߘ�V��:�]m�8B�y.~Sl[[ͱ�(B�K��Co%לJ�J���qԶ��JJM��1�-��<��%M�ռ��6ۅ��m���6�1�q-��6�����uĒ�R��t�۫Cn!�uj<�q�����<m�:�^S�q�q�:�����]~q�!*uq�6y�1Ԭ���J��P�c�q�hqn$␴:��m�q�-jm���%N<��Sd1�N��j�Co!+m���ۮ<�m��!�.���B�Z���� ���1kc�Z^o\J������_�G������\ֿ�-��ο�6�GTK�u�ԅ�J�R�q�)ԥ���:�Θ�����!�:�!����KSKh<��b�SiS�un)J[�)Җ<��u�)jZ�u-�n[m��-n)�q�Jq��X�\B؇��m
Y��ډp�y�ck ۄ%Kc�)�m-��6�ؔ�ՠ�BS�,�Z�b�ZR��[m���۩K�Ω.6�y�㭼�ǒ��R�X�R�(�JK�[d6�:���<��y�R����p�R跛BP�I(y/-�R\ckC�8�m�-��%%�akK�CiSm�����N������cm���yIc�J�q���K�cS�q����-.���K�mKc�S�u(K�l�y��SS�[�[�u��c�S�K�yx�)iB���b�y�J�a[m��T����[ku��c�1���8��a����:�%L?-m���Є�I�?,`ui���97h6aO3N�M�l�䛸cJr-4�sx5Cf#���ݢك��̰�5�-J4�J_!:��kZ�m^JBc�-�1#fTݕiݍ�7riV�W>6u�ԢB�Z��5�R�Bԅ$�	B�alkvK��Kf$�ɳeX��ƼRF����B>u�%�>)kh>BG��)M5j]H)� %�B�Cmj,;��ͧS���E�.�&�M�iX�5����݉c�J~c��ZT����q+CQ��݄�	ÛTي�;�l�Co1�㭿8��I[g�!o<�q����ߛy,c�lyh[����B���b[s\om��Iu�)��-lm	[�m��5�RZ��-�_!�CZJ�SĶaH5hh�<���j�sb���)щ��2�#��Ռc�IR�5YJZP��j!%-iZ��(R���S����)F�F���H<ZQ�mH����k�k_:��%����Xa�ݤ�n�d���i��-ݚ[�a�ճb�1� ��|yLB6�]A�CGPuĵhim$�O�I�Bu-kT��ξK�B�Ƙ��8�����Kf*��ٲ��cv)(8%"�֥��甥!n&Uvh�X�Q���Sf+�L���M��b]��Ɏ�n����~|��u�K�%��y�][jC�6��:�Kq�Є�)y���ևP�{�d8mաkR֤��P��)J��%	R�BT��%))ZФ�*BT�Z��	-JB���hJе�%	��[�$�!MZԵ-)R	IiZ�YhBP��YR���hB��%B�Y(BP�%�iRTB�RJ�������%IJ�vH���B�1Iy
S�	C���)kI&-IBR��D/�1%hBV�)	Bֵ�AB��!*B��������bV�X�͈���M0�X��Z?�ġ5�%H4�	A���RR��Z�֛A���Z��kKu#f��f�c+��5�e�B�<���bZԡ�j��-R\�5VXn���c��M���5(h��6��-,kh�����ٲ��ъi��&���195-KO?%�@�b8�%O1L%La�Ѣl��ѣ�L-�p��݊tulع2Zck&��w;�$��Zֵ-k!IZV�%+R��ku�)+JًCF�/PK�k�)��!��ݱ���lmSvtiM�]ݛ4�ũ�1��j��uš�Z�C�6��C��V��\K�m-���y�8�\~Kͺ���8���!.�HBҔ�եo�m���J�'�l��#Z��R��M���4��x�&���i�N�lv[8\��f�)�9�h:,n����
�ѥ�û��u6i��t����i���M0?>KT��IK]I-i?>m[���#��LWT�iÛF�1�wwl�Lb���ųE�!�P�)|��	QiYIBִ!D,�Є-hZR����`vwilʜ�4�0��Դ5	55�4�kGξK���7p�1N��ɦ��]X�0�ii(֎���ŠKG8��!+B�ƴ�:���&����y��8�l?8��o)�C�<��O%�����1M������[u�T��[~8����u�R�!�BR�����),J҅�1�i6�$��ֶ�Z�ӯ)Mi?�%�%|%��I��8�t���l�)�L<��ZyԴR�����J�Ƙ���j���R�N�m�)���F�X٤�5�:�-�Z�J��$�	ZZ�-�Z�թ�Lc�6cw5ɊwhҘÇWF�N�A�BНm��t���!��ijC���S�IKmR��ԥ�Ku�>JV�)��5�V�i�$�KC���-Cϖ�J1JC�~~~m�1�u�1,u�1*[o�qm(|��c��1��]y�q�y�6�T�1����0�Ķ�C�<�o���z�1�8�-�����!��-	u�)�����u(����KJZ�%B��b�J��%Jbb<�!���c�a�yJB�|���yL�Bu�)��!�����Z_:��h[km.�Z�qM�B��J�V��q��q�� �:ژ��JTJ%,u*C��%/�%�|�P��Yoϔ�:����}�)��c�u.8����mk6�������/-��Qim�)�~S��Z�C��y����������ZԄ��Բ�B�-k%D���D�m(��kRZ��!�jJT���
JP�R�ҢԄ)J-,��+Jҥ%%�hB�BB������L!
J֔%!KZ�B��������R�J������R!Ma���kqhR�SRI�,R�q�����6�B���KZХ$��JP��I+-	J�Z��<��五��)��-$�!���P�
1��y���)Hy�T�8���)�-��>R�� �ZIu�)�6��>JҔ!�ĵ�����b�وS�%�u��!��il�I'��8����%�֤-���K8�ť)YB���iB��%
J�Jҵ!��HcR��)N6�!�O��1)�!O��y�JR�C�$��ی|Kc��C�p�R���_�C�X���chm	Z�ǝq�!����C���d��bV�n����b��8u�C��!"�|�1)u�|ե��~K���!�$�Iq�%oϔ�<����:�-+m�ZB_%-��>|�8jZ��%IY��qHR�c��)ט��C��)�KmN��Q�Ї�BVKV��i)KZ���J��J!%�YH[n?>R�:�P��B��^R����J�ZP�!��<ꐖ��)Jc�)����_-.�Z^R�my$��ꑮ�Ŕ��BR�O�~m�ۨq��q.�jSjS�R�<���6��<뎼S��Կ) �<����+ B�<�K�,�8�V�ԝq�<�<�!�o��-[m�ڜ~KuJC�N�%�%�6�� ��C���A��H|��n�kZ�B:ԥ���hQJR�JP�е �)IYiR\B>A(ZIF�>q���hZ��p��m�>xQLqJ[��$��P�ǜZ�����!,jc�)�.>|��qj[m�ZR�'��ZN�(ZI1�κ�!Iy�6Koϛ|�<�1n5�1�)(|���?8���)�%f�RR�P�-��y��ͭ�m(~Ki?:���!y�%�b^y*q�Ķ㯝qHm/%	J���>i'��)O<�8��$��BTB֤�kR�RP��KRԄ$���-Z�l�I.6�!�i
CR���_%�T����y�BX۪R�	B��hjKK�o>~RT���q/��1�:j�y)q�ڍZѯ��-�8B��:!�|��Ē��JlI�)
~|�%jZ��|��yS���ϔ�!������'�G?���b� �RJű/�BX����д8������n���A�6��ۊ[ku䥨m�Ŷ�%�<��u:�)iq�$����y��!�<�-�/�m�)Ǜmd�ġ���P��m�y���6�6��,S�����!.~m��c�cly�)�K�R~q�-.����͛�V�����bN)ǟ�:���ǔ�o�!�O��u�6��.��JX��SjC�[K�8�<�
qݸ�yָ�☄1q�c�S�l��Ԝy��R��Ŷ�m,1*ChA��[6��8�p��a�m�Iź�CR�)�yn���n��XV�/-�ۋCh:��(Z�6�[�-�B��R�T�͘��E�޼���!LY�J����Ԕ)-���%�j��yM�׈ug�m*Qoͩ����K�ϵ���ל~�%N�iB�~JP�K,�-JZ�JPJ�V��)$�)JR��!KRT�)JR�-Z����Y+AMRP�)%)JIJ��R�%+R֥%I-)JT���IZ��D�d)IJ�)i)D�)ZВ�����!jRֵ!R���R�R�աJRP��d��ڄ-+Bд!IRе�mR�%)ZR�-+J�RJj���HZ�%IR��kZԄ�R�-hRԴ����IJ֥�H)hB�ҕ�� ���-*BҶ���,�!iJ�J��-*R�թ)J��Ҥ��JR��JYJ[�c
ZIB�ĭ+Z��!MJ
R�JR��*A	%
JR��)IhQ-IJZ�R�� ��BV���!)BT�)KB��5(JЕ	R��J�JR�%I-jZZХ��)HR��ֵ�!kJ�J��-IIhZ
IHBTBV�iZ�R�Ք�)!HQ-*%
JRZR�,��IYmB���)jB�(�,�-KR�R�Є�%,�!+ST��
A+BZ��)MJ���BKZе,�Rֲ��%iKP���$��D ��)*Z�����J	QH!*%Z�JԴ�(J�5KJւP-$��QD!
B֔���kZ��KQJR�K���!JZV���)h%)�JV��-R��е%)B�Z�JԔ%(YJZ�AK%R
,�$���,����JJ����zx�Uj����6��%Lb�6�奌q��jq���m��y��-��q�-*[�q'Tġ	B�K�uo!�6��[m���e�!�YL<��:�έ�:�)�<��y�y�1�<�!/)�)�-��o-G�-����N1�%խ��Hu��^cS�cΥn8�5���!Kiǔ����%��إtږ��m��V�K�:�[%�Kq��mjq�l��<b�u-��0�8ym��1èm��-hK�!�a+yD��\c�)���1š�c�K������qKu�֧]R�ŵť�m�����cCBЅ�g\y�V��<yN��q�B�R�ZuM��(����lۮ<�8��\q�<���b�㎺�)��J�a�}M�U~~K�R	mI	R�(��Ԥ$�%IR҆�d-e%+JKRTR�RЄ�jJ��-kJ�-IBP����B���(J�����d�	B��)
J�ZPRVQIJд��)hYY+RP���![�����J!$�K)	R֤�-���1�!KbڂR�$�)HK��i8�PB��-H!1
k�B��	JT��*-IJV�-jR�(@�V��KQ��)N�\B���?�i~JVq�R��-�ߟ)O�� �J�JI/ϔ�VKu)R�JP�:��!��ҟ1jy�)��>R[|��ղ�y�CT�!*u����	1��C��B֦>qJxmŭ|��bT��q�)֤��KZKR��IIZD��	b��B��!(��S5i|�!��>K���Ԥ�|�R�JХQ�_%M�>%���6Ꮫyť�Cn!+S�ІuOm<������%�!n��6��d)kK�c�Tl�(R�%��8�!��T��P�5�u��)򐴸���bԶ�$�>R�����i|�RT���+H��lC�J��:��:��|�P��е��ϔ�?!!��P�!�K�)O�ӫq�)IJP�RҤ�D)KR҂���!e�e�R����җ�xյo<�!o�u����!)�Z�ľB��T��Z�󏔔�c�T�1�)hc��!����-��ZLq�|��y�m�8ĭ�B�J������6�����X�R�))bP��1*bؖ�S[Jַ�	B!.���[m� S_!hm�)��6Z[�R��|y���>BP�Rb��JC�J<���ϔ�%�x��I	R�(��mKP�iRP�-+RR�u)u�-oϔ�R�+JS��J��P��)~|�E��%~R��m�I�b\q�R�j�m���R҄���CZ����
J�Zѯ�|���c�K��RJ_-J�-��K�O������u��ٴ:��E��y�_�y�xšM��f>��Җ�$��|�6ĭ�Sm6�Х8�1*y���q��1jZߘ�6�:�O�Ԕ�V��%yJCc���u(6�)()K R�R�!kY%-�[kS�!kZ���)��HC�<֩�C��!�yB�m����Y�C�V��,S�Z�Z_>8��jS%:�	B��$�V��JZ^B������--���V���ԧ����E?!(c�������Υ��B��╦%�$��ciB[jy+~<�6�ЗV�%�����%�ͺ�%����C�}�!h8R�K�-JP���$��(�ccTBjД�D$�B�ZR�	J��*Z��%D�
R�-D ��KJ�T�$�%
BV�-hZ��-E��JI+%*!!�
B��,���%%������%kJVY+Cy��|�~JB��:�?��bP�!�Bm*BB��)~xRJ%+)*Z��JRԢP�-d-J�ykbԖ-k[;?���!�%[�甦>|��)(C��K�K�ԧ�R��4��<��R��JBB[mJ[μ"�|��/�-HC��K��c�i疷\R�Ju�5-��!�K�m�y
RV�h|���mjC��)M�Ϟb�Z�T��!e�hCR�5+RP�V�����Ї�J�%��o�!�%IC��u��IK����qhyԱq�����~|�K����?-;[���-,q*6��p��k�~K��F��I-�M�lRR�J	C�c����ה�)HC�C椤-���8B����S�q
Q��[�R�����m.��hm�焾RԄ8��I%���և��!*yiB�)�%�"�!�[�n��!��|�����B�K-kI+J	R҅�+-�J��%M���m�(u$�V���xRX�ϞJ�B��1����CI[n+JB!,Jԣm�S:��!m�>BP�|�]x�V��)+Cύ�È|��y��uHq�8�8�t�JR�\t�/�}�����|��u$�����-�mhZ��Z�B���ڌq���S�甧_����kRY��k�
S�%��ͩM���u���_���.8��~RB�Z�|�!!(q0ձ�S�|R�!+Qe!)!
Bҕ�DBR�Ե�%II�ϔ�6�5�Z�|�湬S�R�����J�m��|�<�PĒ�ͭԘu���!/%(b?)Hq.��Z�yJm/�q�Jyn-��!*C�K��L%���,b�ۯ6��|�>C���� �����R��y���~m�������lyĥ�%����M�p�RT��Ĵ�n>R����P��!lm�J|�X��u�ІД!HK��<�(��R�(��KQKR���ZP�KZ�b��C�%ԭ���-iiiB�R���:YKb�4��$�|�!�%�	~|��C�R�ێ%�R�T�����K򍔖1
|�8R�lא>|�-.�H[jS�Է��u�~BV�hZqǟ-hY���T�j�J5ג�j?8����ߊ|�T�<���o���c
J�m���е�~J�JT�??%��~J\R��T� �������hZZ����hJ��iBJ�)IJ�AHJ���%+Zڄ)�� šF����
-
J��ZҒ	AmRZ�T������*B�ZԵ�R��k)hj�Z��)*I-Y+!i%	Zе-�?����RmkZԣ��H~I/䱴6��S���-q/�%
-jRJj֢�P�)JR�Z֔,��-�B�����R��R��ƧP��ה�6|��%IyjChq/:�F-:�!�4�%n-m��|���-kS�R�ڔ�R�M���l�8�\6c��Z[m搗�JꔇͩIj��.��|��Z���|�P�KQO�)Hu	^��~�Pא��[|�R�Ҵ-j%+-	!JJP���,����(Z����[C䥵�O>S��aH~BP���Rĩ)F���Ru�!.)+K�����ڔ�m���mO���y�1�R�^q�<���Д���x�P����(u��K�X�)kZ�m*bV�$��1�J[[�I�ZV��f���K��RcR�:��%�k[m�>R��O�J�Ē�Ÿ�|R��6�%��)Hu)[�)����R<�ה�����8�^k\qkq���Z��Rq���^B��%�!(��jZ����BV�!F)JJ�!n�>R�mJC�'�P-
b�|��ԥ�KRm����*u�3V�䶦�Z�C���!����[�$�I#I�����^yj>y�q/%��q���u��V�-~yî�����!*-�Ty�K[�y.�SkB���O6��~m�Oθ����\~[��u-ԸB�RV�BV�q�-�-�mN��8�����[R^p��N:qM�N5F�ǘ�(�u����Z��PǞShm�8�R���:Ⓐ��ju�X��yM�O�-�P[�~q)c����ߘ��q,mN!ib^yא�!���.:[�[kKB�~m���5�҇��q�!ן������\Z�ſ-�C�S[�.<��Զ�Y�6R�mIZ�<�JR�<��m�Km�Kg�1�(I/���-	[�:�����:��c����\m�Rڔ�-M��KjC�m�lZ�q	[�b���
!�%Ԑ��u-��)-�����6KJ��C��!o�6�1դ�-�^y�)���f�C��{����w��9�hſ?�K�C��?%��[ylYO)�B֦%.���!���y�)k�:�!�R��uHy��Pٷ�c�-�).1m�)%�qO6�qn%IJ����Kt��S�qiC���c��y��:�-�<��8�V[۪y-���!���)�mO6��q�8�l6�-b^[iy���N���p��m�Jc�0��c�b��-kJM��:�[�Z��-��ĸ���)�X���]QG1�-�[o1�8�ż�%jq(Si!u-��[A������!e8��Z�6�yN8�y�J��6���[u�,�M���V�V��ۨuHq()�-n%�:�<��[�0�6��1�)�6�^J[u�:�lbؤ:��-ג��c,��!�u�y�R�Bԗ��1�p�:��]mm��\Cg�|�c�?)N!-ib��d
mS�lZ�bP��b���P���:C�6�8�e6���)
�j�jS��8�!��-jBPê|t�����廬~j�B���)�Km|��uZ�-kST���V��*)k!HR�-(Jִ-8��6����M!
y��|␗��1�yj~AV�o%/�R�~R�>�>AKG>S�S�š�<�X㥭!�S�Z�)�B�|��jc�����R���K�_5����p�ũ�_��n<�n�GXىx��y�͘��b�)Jb�b;*!��o�[B^mjc�%
uQqD�!�b��)LZVK�9��<K��m�Z�hy	C�^�6�X!�)yjS�C��$��%KJT�)+KV��J��)))d)jB�ZT�Ї�J�t�����!�(m�亗�jm�>x$�%�-oϔ�җ����1�����)Hm	t!,~R��R��8�j%��kh|��/��!�%
I*m������B�ZKC���6�E�m,qJsO)H~��S�Ic�-��ϭ��m������_�I+m��/)��l�)y�%D�!IQiB��-$��JjP�)+R�)�Rԅ-*ZԴ!+RZT��� �-k%��%IY(J�ZR��!)J���D)I!+Id)�-jQKBT���)JZ�Z�jPZ��E��)mJII%%���
IK[�J_6~BJT���Z��6�6�%i1HJ[uK-m�q�8A��$�)i%kR��kBR�)J�$������?�)��H|�5�ijS�Z��_>u(Jж>uN�mթ|��ia�4��>y�?)H[m���n)���D��-h|��,��֒��R����S��LlS�%>q(y�Ԇ�C�o�lS��)~BP�R���Z�Rе-kZR���
BVխiJR���
Qd��ߟ)M��-�O<��RR��Ω��[m�>R�պ�1�M��塴��/�~m�1嬗�c
:Kn5�6��q�1�R�~%ԡ-��
u,m+J�)H!D5Ϙ�XԺ���R_�K��|[_�Z��R�V�!�u�JC��T�/��<��X���mO-�Zy֔Q��-/��KR���)�)�jco����Z���b�ķ�R߱#�Θ�:�!JJ��-RЄ!mZҕ�
jP����������	B�R��o�:ڔ�/�y+Z��1|��B��!/ϔ�:��S�jm�S�B��h|���)��>q�P��6�_�cC���?k�y)mz�m���1���<���Kd:����1kBԔ�hAH~B�Jئֳ$�N���yHB����ǐ����[KD���V�Pڒ������%��Z֦�~|�!��5��C�Iy�)֘�V�_�Q*B�(�KJҵ%JBR��d$��+B�k�R��R�o@�!甤?6�:�䡴!�:��B�uJC�%yM�(jKB\)��JP��|�8┄>BP�����RV�6��5/��:ژ����*@۩>S�<�-�)	Ґ�n6Co�C�q��ymt�i~[��m�6�����b[���)C�%�1����Ŷ�<��)��ŭb��>k�i&�N�>R���Ppƺ��Ԥ�,�)�R��-d�e(�!gJ�a�Z�:R����M�C�<������KR~|���b�BP�Ԧ%亵���|�%im�)HC�x�V��J�S��|��1��/�R��R����hRǔ�%��|�)�kChq���i�X�1	b]mjB�Cm�<�X����q��<�%lq�|��!�ǐ�8����P���qn:���ߏk�-)iB���!	I+Z
J��J���*R��HRԢ���k,�!kZT���%D�SP��iAJRԤ��ԕ�+Rҵ)*Rҥ-JB�BT!ZB�IhR�)IZҒJB���B�JҢД!IZV�����)�o�BBڐ�X��e��ZV���6�)o�8^��iRP�P��jBT��JB��(���-H~-hZԖ�:��jR�ơHbT�?:m��iJ[m��Dj�V���R�T�m1��|���Jb��������C�J1�ҧ��%��tQ���T���R8%(~BP��8ĥ(A�>|��1�u	ZX�JZ^RT��|��-iJ��)JB�)JJ�QJ��KK	K��>R��P�-/4��ה�>Z�V�!����N������o?6�<�c�%O!�疅?)�Ÿ��][�����5n�)*~C��)
 �Bև䤤����%�8�N��R��)��)��R��:��-ġ�<�V└5/�����8K��R���Z�:�ju�)�qHi,Q*|��Ω%��N�!(SN�kB�)LyJcZ��Ї���jB��%(Ae���BV����
bօ1�J�_>yk|Լ�!�����)����(�6���JC�+\5hS��җ͖�$��|�!�K��ο:��Z��1�[�_mH|�-,-��8�c�O:ĭn)	~[q��f�8�ͺ��KP�F�j�X�ԧCi ����0�6���yLե�J��<�е��kl���>~m�y$�BXk�-o��	p���3H|┇��S)Ly�hԤ�i6|[��IY+RZ����+JҕZ֔��-ձLRΡ!,qJC�<j��T�R_�)亥-jc���-H|�P�M�K�u�Д���	u+ukJԭ����#_!��-jZ�:��RTJ�%��ֽb[u�!�|���!�XuN:�n�ն�n�BY�8�o6��bP������mz��6qM�d��)hj��%J�KKV�!�?!��%�8�--��R��n-o�)Hy$����<��)*BTS椂�-J!e-�RP�Ql-(B��)��R_1O�Z^J]p��P�%���J~J^Q*J�������>a��IR���R��^k�_-O<�!��q��J[BxBD<�����/����%��:K󏒔��)O4�]Z���%Z�Oh�)Կ)ImLI��S��)��S�[�m	8��������\Cd-Ժ�m��m��R�T�o���X����QHy���[��ҵ8Ǜqm����y�)LC�<�qE)��iqM��έ��6������o�-g]qŭ�Ē�-M����k[���]c�[�y֧�S�q�:�����q�?%��\y��Y��)N�q�qԥFҔ1�LY��<�V�n8�m�ۨS�6�V��Z��Rm�8�6�iB�6ڝZ�yiu�)	cJ^@�Ҧж8�XS����)n�����mǈ%n!��y�Ժ���C�R�y�%iZPזŒ���m/�c��ߝJ�8���q�1�6���RR�(�1u
b�Q.S�Τ�Ԗ-�V�V�%n�8�š������8�ka�6�%䘧�8ǐ�ha�T��?:��m�8�?:�!�矧�z�)�S�%B��:�)�%hJ��KB���hJKB���!BЕBԥ!jYjJ�Z҅-JZԔ�Zҵ��)HBT��J)�Z
%e�JIiR�Zօ�-A	Qd!KQjJR� ��	R�JT�)+jR�,�աhA*BT��	JФ�(RR��
Bҥ���iJ��P������֥-KJT����R���)JII%$!�R�Rԅ�*B��!IjR��R�$��)�BRV���%JIh)J!�Z�J�P����%�+JRQkR�յjIhZ���BHRЅ)KZ�B�!IBT��+[R��h%jY$�Ц�B�� ��R���
SP��(QiB֥�j���%J,��ZT��hB�Z�J҄�(!Zք���+-*R�JT���V������iR҅%*)kCR��IRV�)Zҵ)KAZ��Rڤ�Q+J�CR�)
JIB�R�������e�������	-jKTZI%e�*ZT�!�ZЄ!D�� ����
R��Z��jjԔ%J֖��-�JZ�Ik%KZԢ��%*BR�!D,��(J��!+ZR�%(%KR��MZ���-)J�)E-�JTQkKV�����+)
RT��
QD-j-�!kj�j�%IR�5KAQ
A)kZ���-JZ����-+)*J�ZĖ�%+B���l�g�F:�)+|�>m)O8�-n����]m�qM��_:���%�P���X�뎼�l��c�u���1�1���ļJ�B��ĺ���l)c��qmS�]y��\B[�8y��t�Cyԡא�ж<�R�m.�
[��bq�<�(�um���S��ڊu�m�ZЇ��%�\a�ִ6ꘄ��:�:��BuŸ�V�����M��C��yn��j\u嬇P�\yM��q%�N-�����bв����<�n����-�Skc���jBu��q���m)c�JT��N�<��q��a�-o!m��c��ylc�y�!�Z�ǒ��כm�[l�Ckm����)�Y��Os_qh[�B��k-Bҕ-)B���*BV�AhJKT�)E-KR���$��*Q*R��ԡ
-�%�(B��5kJ�)jP�!J-mQ-J[V�-�Z�IZ��!iB��!j!*Bҕ$�ҒVԨ�T���V�إQҒ�)�6��␇Z�d!c�)uBKR�J҅�	I)ZTJԵ!IB�-HZP����8�)��B��R�:�)�kB��<��%hChJߟ-kK�R�A���ҷ[C䥌R�[�iOϛR���y�jJVR�ԏ�buN(�>Z��I<�����hR�oϔ�?5H|��b����_CTuC����A(-(R��!RT����*CmKYLRVb�R�ĺ�>Q��<�!>u��򖵡������J��<�!����m(%�Ķ�6�:������Μb����!����8�!hy��+-/�q�~qKKiR
R��T�!hR�6���ku%�ͩZ�Rԡ�/ϐ�T����)M��:��E)���hK�C�|��n��%��JqJC䶤8��mKC��<��HJ��>BP��bЗ�R�I(l|�����Ք�-kJT�)JZT�V�,�(�)RԖ-KC�R�ԧ��~jڔ<��)[��!iB�ߟ-Mj�J6�!�����j-�YM�yHB[m��:�<ㄩ�)���A/�S��m�T���-�Z�[�u���C��q򐤿6��~8�N-���LC�1kS���uHZ���)�j!ӋY�����RJV�Jlu��:��І��^B���-���m��!�)Hm�j:~aG�B�)IR����-iJ�)	Jԅ-hj��))�_)N8�!��H'T�$��|��uHZP㏒K��-Sn�HZR��٫j_>qykZ�!����k��Ԓ��Ͷ�<���n��)+mJ~|�3O6�:�?1�_�-���Ͷ�P�m�-I����!�n<��yO�<�V�:������BP�M�HB��1�c�-~KR�X�(�)���T�փ�7��k�_��!n!琅�?k�R�C�%~R��e)�����5��!SP�-HjPRԥ$��ikhb��)Rq���R��%�P��<򔏐|�O)+1Ժ�k5ZJT��[�)N�ԵJ%��<�����!�R�]R����>BзT�?%����Lt���k[�-H|�X$�?�_8���(Km�_(�<אSK�)S�S
m�_���>u�6�ĥLu���mO�q�C��uhuo:��!h~|�8��5	!�S�%+)HY%E-Q+RT�-+Z��%IR֕�IRV�-(B�J�Z�����K[PJV�-jQkR�֥�JP��hR���kJV�KK)+Id�����+Y(ZT��K%+B�I*J�J���������?)h1n)�mN�|�k1t���,R���!m�!�/��䐕�����Z��!
R�B��	R���	S�IwR�!*u�Q�C�%ϜKέ([m��ĊCR��)Hy%���k���bR� �ߟ-Kk�'L-(#Z���:��0��K���1KJ]BP��
P���-o��xꖳ��QЃh[��[k�k�>yJHYe�i-JRJR���(Akq�K�)�bq�į_!橧[IN���&�|��!��Ԥ%��~y��ϒ�j~C�qy�<�P���؇T�6��lZ���Ї璔)y/��1h1(B��/�J��m�N-'yh~j�u��ZP��q�uhi->CK4��d%�Lӧ�ԏ�m��m/�5-<�V�o�JV���3P��JS��yY�Q��lA	BVI(!D�%)
RҔ�JII%Ɣ�!l-(S>KlK�1JJ���A�ZҌ|�/ q~Z^y���>|�)Kc�1.1玶���6�C�u.!�m)q�:���/�~[n�/�?<���)���ļ�%�YHYN%HbJQN!(m�P��!��P����u�!�P��m�%5���)�Ҷ%�5�$�ۯ��K[u�@��ľAhS�Q���KV�!+J�hX�-j!
%-�kJX��8�.�ڏ�b��.>|�T�iC��Oơ��1Ծq*u.4�>q/�S�R�>B�K���iGϒ�����%(Cj�M���[Z[�:�	S�-�S�_1n�q�hf��6�����m���q*m���)-u��)�Bڤ��J
b�;mo6�lZ�8űh-(iJy��b	j��6��KũM�����i�5O��-���hkĺJ��RҴ%*!jRPJ�J�8�!
,ĩ��>Q�)�k^y.>|p��f��x�R�>K���q��!)Zu�V�%��-[�S����N>S�����j�K��|�<��,|����!F�J���Ը�-�����
c�8��S�V��m�<�`�u/5���K�%+K�RC��K]J�-(JP��*Y
B�����Q
JV����I%HJ�ZZ�B��e�h,��%(AkA*YK,��iB���5	)iZ���ZJR�-	Y�J� ����e(���Q*JHQ
Bе�	R��)+YR�c�pR��N?!bP�-�!�b��-jb�mhCT�ԅ8Sd�m�ib���IBP�)	JRRխjB��!-	miR�%h[C�Jؗ��)����u��ZT�1�$�ԧ��<��CT�1�+ZX��/��TJ^Jhm�S���lꖶ8|�&��Ia�y仮�����Z�y��sVKIB�KΤ����AH[TB�Ք��+B�QJBօ�SmJVc����uN6���4�J�byKn>J�~x��|��S��1��V��JIx�ք���Oͺ|����RC��l�����KAh8�jB�!([m��X�m���Z�Y(iŤ�����hK��i���T�	c�5M�҇�S�m���RT�R�Z�����>Kn�%�k���a/��J:�y%5�%��:��ij����O�R��K �ЂV�-HJ�B
Cj-lJJX���)���6��mu�!q	[<�a������~1Ju����!��u5\ޢv�H|꒧ϛ|� ��CK��@���C�?<�c��u�I���_�b����)����Ciq/:�طC��6�8�X��Z�%�8��S�m�1�6�m�z�ڥ���[C�1���<�8�X���[gZ]y�S�:�n�(S����cέM�)C�8�1:�J[b�cX�R�8�%,~BX���O?8�����R��z�)LcN�甅%�~%.�j��C����:�%ly�!,Y!���6ۋZI-��[�!ŭ��b�q��S�l�!.�IRۍ��TJ�[�8�8�y�u.!�)�:�ص6����S�%�)��8�Co$�<b�Xǎ-�q���y�Iq-O-�yIu)y.-/:��1K)M�ż��c�y�<㮩m�Լ��8���5�lu�T���%����֣�c�m�5�91�)o�!��C�:��uO0���,��m��M��m�R��q�:�b�[Ω,ulc�I/1�1/%ly�J�q�-���Z�ڜQ-�.0�n5�%Ĩ�םB�Bu�yG��T��C�J\m�[�Z�m<�\b���q,B�ClSͩkl�mhyfֆ �:�q�)�m��V���Iu�:��[���m�%iulyLyn)Ǜy���<�8���Kug:��X��:�R�Y��)%8�6�y$�fmז��)!�<�1�1�)כuD6�T�V[�8����J�BZǐĶ�ڒp����Lqה�y�)i6u/1�ZP�ic�B��X�n��l���ǜZ�S�B�ĭǝ<�X�^q�ZӮ��<��BԒ�ĞCh,�!d5ԥ���ChbZHB��!	%BP��1/�1�j����O�q�P��|�%�����_:�q�,��%����j]Z_�|��Є:�5JQ�
JR����%jB����-	S�1��7�bR����k�S��%�J֖k_<F��Zt��'���5!�o8ڐ�),|�[����4��~IhK�-�R���5�O�q?%�6��bN:��C�䭷��
kź�V�C��b����Ԕ����=���T��e1�8���	RPԸ��-+[���!�m%1-bR�T�BA�8��C�д�/�Ͷ��
B�+R�V���-�?$�RԝC�%���qk��[�-��-,Z�)d�%��-%��-�[4IR�!kA��m
�:�X�?8��J���<|��-:�X�]m�!�(K4��ۊSZ�>B�K�Ρ���!lu�5��[i|�?!%���!��:�)��x��Zu�[了��!�P��o�[�6�6���:�<��6򵭾J�?8����^$��P�:�-I[V��+!K)
J�-jZZVԩ*ZP�-iJ�-j%E)(JR��B�SPR��!jAZ҅,�%e)jT�B�JI!d�kR������KZ� �е�(�����	J�!)B�������(jЧϐ�-IJ�~[�!g���o!�-��~bG�u!��q-Z1�)iB������LCo-�~RJ�)JZ�����%(Y((�0��	!��,K��|k�i!�?8�_�����K�4�y��[Z���0�Z���'p��c�lS�ϐ���C�CG_��),kPםN����|�)if��Ω����>AO�)����:��>J��KA%��I!�mB��HQ��1�ԣ\qI�>x$y�m�����0�y�~K�-�P��C�:��y����X�m�]J��[m�:��C�mM~S��<���W��]~y�R�Z�~SR���1ĵHm	R��1�5�R(�!Hk�Y!+u6�5�%E5�4��V�ԗ�5�>C��IZ������iQ�i��O ��X|��Jc���i|��ΠH��͞u�iB�|���PAo��ƟR[|�!+)J�Bֲ�Z���)jBV�[5zZ�J����N!�~A�5��.����KZ��^5mihK�)�RèjZ~y������K�K�m)�u����:��/8��y��R�X��ly�1�
ZmlY�BHc��[��O�B��qn!���[~ck0��h)�-ŋJR��6�R��1��Z�IJi��m���A��|��~~?%	m��H���I�6 �V�~|K�Yl>A�Ж�m/���Ʃ|�)BP��J�ԩh-�)KA%hR��b�1*S�mI~|�5� ����	c���lK��ֺ��R|�iy(JX��:��KA-?).���CiR��@��m	|�:պ�:���~J%���p����~m
JV��)ǒ�?)š�_:�д�(��Ҳ�JZİۤ��%K��+B�q�YhKiZ�Z\[|�V��^B؄:�Υ���icQNC��B:��(IKR�R��!�ZR��JBTq���b�8ۯ�)���B�y-)�KjS��l��Y��Kn�:��!/>kkq-H��������)��B����)KBX�P����>Km!��~[��-J���bZ�RT��FБ��c�<Đ������U!.���8��T���Y�5Լ�<QJ!�[T���)(R�%HRֲ���YE%e�I-*!+AiJV��-iJ�QKRJZ�!�R�J�Zԕ�E-jBPB֥��)J҅���$!ISP�����R!)Rք�jJ�AkJ�R���%E���I(��!�)�O��b���b�8�ւ�J�RPaC�-��o�)���6��X��	<�1HJ��iJT����	Y*BJYhC��e���>~uG�>b��%�Cmk�8cn!.�Kc��x@u��^Kbp�ϐ�Bփ��m��b\y,C��]-,m�4���O�شֺ��c���K|�wRjI�4���h6��$��(J��)i)d-+R҄�HB�IjC���%lZ� ���ֵ&�b_>C琧T�0��?$�Ї��矟-���q�^ciq���o�J^~q���y����u)!�������5*y
6�(���-)KkB���5(��E��|���y�O1	~<BX��i�~�4~|��|�-���!��C_>I��� �PD��!���)	qjcϒy�k\C�%�ۮ�A?(��|�,RХ�jjД���kH)LK
bm�T���Sӆ����ۏ��-,q�m��C^S�ر�����,�Kzq,c�����?-�M�	C��c�S�K�m��kyN<ĩi[��mo�y/�y䱏-��H~AIyiRz|~m�!�͸[jS�Q|���1�$�1-ձ��i$԰�Ԗ�$�8�lBA�%�ߒ��^c�_)�K}��Rֿ ���1�@[�x���IR�j5�^5�ľ|��68����KJ�%MYe��V����kBԔ�!kb�%*c�)iq��)�ĵF����R-L~|��!���C�>mj~J��ְ��җT�1���\u�j���K�'N�|q�-ht����Ժ�>K�κ��ͼ��,qe��>~cd�k��6��_���0��-/���!��JRI	~R[J	BR��)BZ�� �1,ClaLq.���C��B��%��"Co%���m�R��B�RP��%d�%D�iZJR	)n��[K?%�$��5-j�Ko���B���<֠�8��K�cHy��<��L>B�K�!�|�]CR��>R!,pA������-����6��!jS�%�khjߒ��ےk��u����[��ߜB�K^q�!�!� �6����S�!R���.6�V�8���?8���C��cg���)hmi[n��^b�[�j�<��Akum���<�y�8�mm����6ǔ����-N)�T�[c�c��<��Լ���R\�����6����6��-�Hx��뒗V����~qO?~b��^c�p����ClA1�)ku�m�,����CjuO�~~u��q�Ǜp���jSkB��K�<��]S�:��T��R�1N�	y.5�-�m����:ޡ�9�q-Cn!�[�y�8�Ÿ�)�yn��an%q�1)So�q:�[y��<�������m�km!�1m��Z�^R�b�cn�%hJ�Y�[)*uN�c�)jy��][l�o8m.���/%KZ�!�Rb�ZM��%�V�u%���u�)���Kn+��o��n6�RХ�������JQZԕ(��R֒�)I!B�Z���e �,��jZV���+%Q*IJRR��%-B��������R��%+BԢ��)+B��-jZBR��kJ��խ)ZR�R��)JJ�)E��Ԣ�A$��I(KT�����-Jд%+)jB��������J
%(JRԔ%kJ�!*jԄ�%(Q�HZV���-)iJ��,��V���$��iB����j!jJB��-hR
!IZ�-K!
Y()d�(JT��YE-%%*R���B����R�Z��-)QZ��!jR���%(JւR�Ҵ���$�jJ��*ZP��kR�%
Q*ZV�%jBZ�(�֢KZ���jZ֥�iZj	RJ���jJ���))ZR�A*J���AE-+J��!�Jе-*B��Ք��J҂�J���(B���YkAiZ���IJ������$����j-H(�ִ-
!iJ��KRԅ)-*Y$�+BЅ���Ѕ!D-D��-hQhJVZ��%(!mY*R�J�����Q(��	)KR�JҔ)jB����d�!*%�I([V��D)$,� ��� ���-BJ��!+B	B�B֤�*jҵ��!E%hBIJP�)K!IZV��B�Rք5
R�ZR�%JJZ� ��kRP��q/:��m*u�u�8���:��y��8���:�!O,�V�(یu�[ͭ�����h6ۄ<�Ω�y�6�<ٷ��8[lRM��R�C��Sm�n8��-����qN��8�6æ�ĸ�㎱�]B�Y,y�C[q�J���o-ա%:�N!.,�n��O:�%�5jJ^S���[�Iԩ�-(S�mטî�J�qLy�ĺ�:��m����[�A�)	q(��u-�mm�Sy�l[ěy����Ku�-���8Š�1��6��qǘJ�C[���%.���u,mKR[J�b�c�B[	u	u.8��mf�u�<���J��<��qN����u�%)!*1����l6�S�6y�-�^q�c�<��8�mo+\ӮRb�KIեkI%�hB�-h)+R���!KRR��)J� �-hJ�-B�-Z	R�YjB���jBT�д��R�RԤ-IJIBR�$�$��k(�R�*R�RЄ ���������-
R�%$�d�+IkB�BP����ͺS�C͊R�a���!�B�c�)�)�kJ�J��]m�1hy.�Jm���[Jխ�RTZ֤�
R-e��PJ����גq���>k��_����6�(Ƹ��m[ZJR��u�~CR���ZX�䱉t����X����Km��֥�q�]bO�؁o%�?%��Ja�5N%�4��5�1�� ��J�J�JšjZ��h,q�RP��(Z��o��C�_$��� �6�)
R�|�q	m��y�8�B��S��0���Ŀ%LmԱ.k���~ycm�u�m�o�%��b[b�,�!	K�p�6��Q��G]u�,�^:�\@c�~~I��H"��C�~0����[Aֵ���<��6�R�����Zy�O!��ƞBZ?):��!�I[[~K���iq�k_6�!�Ρ*RV��kZԅ ��B����iB�h�0�)K|����;���K�����%�8���4qğ!հ�մ��ψykZ�Ko�P������gͬ����~|�?6�']m�c�cS?>ulq$%KZRJTژ�6����-�?8��X�mK�Q�b�\m�<�)�%���b!�R�Ķ�!�|���Ic�ZKFؗ��bJ�O�>m[�e �-hBЄ�JJ֔%)Z�BԵ!m�K����%�j_�~A�!��6�����>K�֐���y���ҏ���k���hu��J���k�|Z��hi�R҃�)N8�!�渄��lBߔ���JϞy�uO)���n,��K��o��5�Iu������4���덥JCq�Ĩ�IIB
J��1�[[c�%-��m�1�?:�:~x�+_�S��]u'�8���Pb��>!O%J)JR��KJRYd�խ&��%lB֖>CV��tԎ1/���:�)(a���V�LK��Cbu��o���L|�).5���y	8���+c�!�ϒq�'L~A-k�4�Z6�%�-���y�h�R�iu�u�/�l��L��RR�-�6������V�����6��B�B[!��	J����)hj֕�k)JJ֕�j!hB֕���iJԅ�
!I-iB�JV�P��$��D�-hB�-(Q	Z��KJ
J��hR�JԵ��ք�+ZT��)RR�֤)kB��!($��,�!D�K-jjڵ$��kuJ?)���-
|a)uHJVK�)k�mkZX���+u�$��jҴ�kj������RV�1�aR��|�N!�ҚםJ���㮩K|�T�O�uL5C^�:��%��6�X�]k�jZ��-kSoωq�icd�8��C8���:�]~8�
yJC5���[�/P�k]Z_>I�!��?A���+!hI
RT�%iB�R�-�X�!ia*C~B[cz���m�4����m�B�K��)OK�u�?>|�Ғ�b���q�屵��:��V�J�C��8�o-Ԓ���-LSk�|��-,b�KkRքJ8�4橦��\B�R�c��8�[�6�^K�ly�P�%�Mk����)A^u'�[p�����K��I��!icO�:��HZR�)	Z�IQJZ�Y*BԵ���ԘY�B����O�5-c5L~q�򖤰��#Mk�>J�J��?<�/KfЦ����y�|��?-iK�uFϟ1���0��m���~%�JZ^Z�����8��8�bХ�[n����� �Tb��JԆ�,Q,[Z�7�Zۭ�qIJT�ߚI���S�����%,-�)+|�.<��u~b_!����Pڝ)IZ���KRҢI*Rօ�
lAkZX�-,~|��ԭ��(<�]!��K�-��m�,֭�.<��?(�|�^RҖ<�X�]ii�4S�[�|��))Km�Ibk���|�)�$���?!���:�X��yM�N:�/_:���G�!�J�� ���┅�Q�1�C�8��)m>AkkZ�q�ΝR����	~|j�N%��X�5��o�JФ$���)	J��%�ZԂ҅���1hSS�����5f�(-��ix�X��kImi*K��m-5oϛJ�-(c��mZ�ϔ�KZ^C����J[B�ֿ>I�iO����^N�~m�R�� ��|�Z<��/:��K�c�ϜRP�ċSoμ��kiu��b�:�s�C�PB��?!�hJ[Jԥ�	,��-IB����*JTZ�!HRҕ)*A)BԄ�
Rҕ)*R�5jJHSPBIB��)K[R���%�Jԅ%$��IB��ZR�%e)HB�B��,�(��kR
JR��+JP�P�!(B���)+BP�!!�mJJ�%�AkS��M�LbR�%+[n%�6�_�a�P�ԅ�jR���e!+Z�)KQ
Z�)�Z��RX���1��!!��|x󥱷)Hk\u'�sV�b�>m��_���,|��nֿ!N%o|��Km��$!�K��q��C]q�%�Jc�::�>KUf��_�%�#I5n���!NJ���)jJHJ��!ikT[�0�������5O�Pג��6꒥��ϒ�ͭ�������6��ז�[��B[B�u+Z���b����θ��Ku/ζ��?)�>S�C͔�K�%�<���CP��m(m(6�6���4�:���_�CZb�x�X�5��m��J|�8�Ο8�V��֘��#_<ީ�R�uZkK>|�?��K�!�kN8�!����lC�]B�K�Z�J�J��(YJZT�!Iq�-lY�Rж>CTľS�ym5uN?:�<�!��8�(Ƶ�Z_�%��$�Z�HB�����X�	bY�~�L)���[��u�kC�C�1�6�k|��uE��<�n!�S�hqm�m��,u%���qOζ���R�{T�Ao�~chZ��6�n���㮼��!.�B��T��m�1��q!�C�B��J^u���1E�8�:�n����R��o)/%�,��ոï�T�R�yN�	t�C���u���~<�<�jK������!��T��6�%��Z�ť���n!)yMB��-/!.�	u*ZѪSY%8�:�1.��1�J��n�8�!�:�����ߛb�y��ſ1,c����:��B�mmM���{R��O8�?)O%n%�?%�X�����[��1lm�إ!��Cf���<�KfاT����[ILc�-�8��C�-�����!kR�~m�5m�S���덥(m&��κ�)+Z�۩qο~�T~y)u�۩[�<�	b\J֢��Ԥ�����jSR�qա�<�6m/-<�X�R�m����hy)�S�:�:۫u��������ם[n(�)+y�:��ujC�8Am�8�B��[������\C�!)k�-/1�m�b�SQn-�8�)Ǐ(���\Bж-Ű�]u�8�Z�y�P��!o1JyC�co<B�!�:���-���m�S�cd��a��%�Z�^y
qJy*cn�ؕ)-��1BP�$�V�uա)ulC�u	m��Ę�:�6�8��c��I[n!�<����u�)d��!O%GT��ŶĠ���c�V�V8۬[m��B]So!HK�q�mB�X�c�1iqI՞%�\p������Rb��)�����%IA
P���6�8፬�1_1��և�BR�1ǐ�������X :����[JZP���jӈS��[@���-t�)MJք)jB�Z��	Z�ԭ)lԱhZTƱ��t�P��Q�q�m�|��,m�� �B��qO��?0j���<�f8�-��ZCMs_'O6�5z|���%KZR��אJ�)��C��ϒ|��wPR[|���꟒��۪~m�8�[C����n-���[iuiS�n8�5	BP�R^m�C�Jm�-N�n6��q�Kkjִ-�)Ic�)�>Z]6��Bè|�8ľ|��6-����JIB҄%�J��������-&���S�T�>BV���x�O!G�_%�?>K� ӈ-�^`I�?>u�1��LtԚu�|ĩ����!.��Cf�!-|�P�0�5��~yE:�:��,|�V���f��KB�bҕ:� ����Kϒ�Ԙq��!�%����iZC�sju���-E���jQ$�JZж���*j�Z�R��!KJ�R���k%BRRJڄ5)!ҥ�JJ��-R֔�d�B�!*Zԅ$�%jR��5	JK%�j�Ԥ�HBւ�B��-JZP�-d�IR����Ж�+~>y���1M�Ky6q��cζî~K�A/6��z�kBR��CRZ��ҥ��R��))K�J��0�>|���I��V�6��亥-ia��ֵ1*|���������<�)�>p��%-%�|�O ���K�RR�8ZZ��1��~J�H���<�R����%�P֎ �i[�ꔤ5����u(BRB�JYD%ij��D����J�S�>|��%�Қk�%��)/�BC�N6BP�E��y甗ĺ�y��8�X��,��q�N8�q�6���K�%��N������Ԣ����BP��|��֟��ZX�V�[i �t��%L|�Xĺ@|���%��Bζ�Pk]|�]I��Hז��μ�Е�>A桭1�|�:�4��:|�J���IJE%h!)Z�! ��b�b����/Ϟ��0���)S���@�Lm-�$�g�Q���)��>u&Ї�X��Cm�%�>m�X�Kc�C�j|�M���yz��|��)R�(�1�<�kb�B��1KR�Si'M����Э-��)KCi5��M�*|�iגq���)
�>u(K�:��k�c��5����դ��������+ZR�҄�Z�6ii1lJҖ8�.6��<��HuIS�?>!�[u�]kPk^םQ��m)�<�Rꖴ�|�jp�>B�J�y��Q,u�$>CK��C����ۏ��|�o:�ϐ�<�庇\uM��1�m�-����[Y��Y�>Cl�8��1��!�(�1���8��J���jcϞm
R��+^|��kZ����X����ԟ>Jԅ�RФ�kI	)K%HI)lj����JR�6�� �L>qJVy�i|��!��K�@KMBJ_6��K�5�_�8�>1>y.:���|��In1��P�1�P<�6��6khk�j�k�%���׋1�_)�Z�If��'�1i~qlCC��m���שRC�-�屍��'��1/α�Jy�y����P�:��PRP��B���D�jJ�B��!	J҅ ��k-+ZХ)I�-KJ��$���%	B���))kZ҂��Ҵ%JV���+B�Jڕ%% ����	ZP�!+B�RKJJV��ICP��)BR�B�%�B��%.�y(J��P�%IjR��BT�q�I�5	m)6�hJR�RR�RT���%Q,�����K�),%8��5-5n�������5�1*~|��cD��8���ԡ*c�:��Q�|��~[�|�6R^�س��cZ|��AţRƐ���~q/�Z�6����48��K�%�P��ϝyn-+b�!KQj%)RP��
B�Z�Y,h�))c� ��-�O??5��$�O�u+JX���yľB�S��^c�y�t��R��J��q�bKlȓ�%䒔��
J��%�y�KjchCiShY
`�ͤ���N�ֿ���_��ix����1�)��<�%HR؆��klS�1�%�{[yM��%
Q,>C�j�sT��/ �k��<��BT��JIh-JCP��)(��B[i�c��iCB����q�F�>co)jR���c�C�k-LH�B�֡�ϝt�)Im��M�m�n!�VQKch8�o�6�-Jmo���<��c�K�1Ķġ�%.��)�O�y��b�m�:��Cm�N �1,[�qK�Rk_-�O�%�N8���� �亄j_)�j<�Lq�ϐ��Lq�S��]B�8�_!�m,ig>R��R֥-�JIZ�Z�Z���ա6kR�����i>x��y/�:K�ġ��x�%����B]Km~C_�CPy���BX~CkK� k�伂����B�6m
CJ5���8��%����ukq,uխ���|mjc�k��6�����_����嘅�����h[�T��ĥN<�u�1Կ1/���-�y*SR�$�8���X���khJ�<�<ZX��_5O�S�y���|��^�����%HR�JV�%e-KRҥ�hR�Z����LR�0���>I�)��4��oP��%n�,k��k�-��]J_%�u�8jk��C�BXۯ��cX�5�
CK~|Cı֐5��~םQ�5�RkX��?%�-[���-�S�:�5HeG�Ω	q%���~u��%M��uk[�:��+m$0�^S�Jm����u*�>S󎡚�ߘ�T�?)�6�!kB��y����$�-l�:�R��yĵO%աǐ����),S�Sv��[���1�ű甤:����b�q���-�[mŭ丵S�ck2�K�%ǌuא��N�[[�<��x��b�KjJP��8�����㎸�[�K�m�Kb�b]Ju*q�1��iu�_��mn��͛y�hy�!�X��[�����]u)Kh1��<�q��q��k8��m/:ǛJ��B��R�=�yԡ	y�<���R��ַ���q����P��:�_�qyJt����1n6�ǘl�T�T���ձ�6�ߒ�[e:�u�8�~K%iz5��cθ��8�ĺ��([�qǞy�CX���<��K��K^S�B�hy$:�Z�Y�!�ZN���~B����{uc�R�%HJ��V�)e���(Z��,��%KZ
)h%)Bж�)Z�,��JZ���jJT��jRT�%)jTZ���hQjIR�-HB�J���������KBBT�!R��-KR�,��%,��Y!A
Z�RP�����IRR�-iJ��
A))IkBBT��%�)Z��(�	R	jV����
J��J!
IkZ���hRJJB�ZЕ����V��h%iJ
ZQkZ�)�IR��)!IRJYiBT�5KR���	BT� JJе!	R��%)-BԴ�D �!*-IJ�ԐJ�Z���I	BҴ-*Z�!Z�(��ICVBֵ%iB�R������!KS_�QHA,(�RP�)%�	KP�)jj��-E�����ZT��	!RP�T����RR� �!)RP!)YhJ���D�KZV���R����IR�Z��HZ���k%HJԂд��5jR���Z�%jBZԅ��!D�* ��
Z�խH��(JH%HQjZԥ�Z�J�����Ԕ5+)d!I�jYD ��*jP�!HZ�Z����ւV��$(�����$���)-h)kA$,�Ҥ��-+R�BT�HJ�RV�(����	I(RJZ�!
Z���JJP�5
B�д��,��+J֔-( ��D)iJ��%+R���KBԴ�z#�[�\B�Ϳ<���<�^mO1�%e!u��K�6��x�m�Zq�8��]J�[n0ĩ������qbZ<�Z���S�m�Ʊĸ�P��.-���!�:�֒c�<ũ*q�]Z��m�lu�%LB�S����:�n6������6yO��<�8��q�0��(��yKΡ�:�uD�lq)J6qk[n��X�κ�Lu��S�u(S�8�mHm-��O1��:⒒t��y+q�hp�0�1i[�[�-n<�1�%O6�n�����!��ujZ�R]B���]uF؇��Iu�1iq�ı�cg�^Sm�C�[!�kAFж-O!��B�Z�p�]q
k�aIuo<��y���]m�ǈcm�՞<�qHS�}�k���~~S����B�B�!I%JB�����!K!HYj!jB���jP�$�)(RTBТ���(Z������)(Y�+JT�)d�IQkJ��!iBԕ�(ZR�5i)$�%)))
RR�,��Jե[P���(B�R��丗�kl[�ԅ��)�-m�8����BT�%�RKR���%	Z���Z�����J)li�ԭ,a)R�N��!m�����Y�y1���ԕ���xޱ�q/����<���A�n%!,~|�]I.�KJ5��K���6�%IK5���)ĭ�V֞y.?6���c\~K�@�!����6�><�R��)AHJ�Z�-$�$��!*84�)hbV��ڵ��ZS�� �E�%���C�Z��%�u,S|�����8�y<��?��S��%�?6���z��طC�!R���J�թ��m��[�T�iqÏ�8��S�qD6�KB_>h���>K�Cġ��KV�ڦ��uiy����)��֟!LK���P%�����?>C�B��P�=�iLK��?!��c��B�-)BT�-)-D)iJ���D)hB�8kP���������8��0�>�䨵�J[)�-�ϒ�i�P��y����ֵ���<��q-�Kq��ϒ|�Lm��KX�6�-��ǝ^��:���<�~b�c�I���َ��1j|�X�����6�8�O�!����>>CRi�%����j�Ը���Z��%��HԺ��%԰��d��+J��%Y	)J��HYD)$��Z�1D-L/R�>CT�_:ԠCZ�Z�y���k[�񨦵�b_���������)Hc�1iq�C�%���;��m�BX�!���/!��K�?:��%�%l|�)��K�:��<S��%O�mN�mLR�����^B�~J	~j_�!�-	|[�!'T�҂д!!+IKA+lֱ�:Sm����l��kP�O���l|�ǝJHB�V��IiZԔ)iZڢJ�kHR�ŭK1�Υ�|��M~,ּ��:�RR�%��$�Aտ!�i��u��jI��K�V��>JV�X��P�� �:kO�mi|ġ��iyE��^��?:���-Ja��P�j��>|�k�}�Cn%+l�(�6��� �q�TS������N)㮶���\��P��p��+YkR��Z�!%�+Bд��KR��KJ����hJ�[T��JJQI%JBZ��)ZP���+Z����(A((�҅!Ij����KZ��BT��II+J�Ԓ�%%���ZԄ�jJV��),���m(|�����ڲ��5RCR�� ����BV��ISV���)hBR��)ZЗZ0�-J�ͼ�ؗ�%�y�>yIp���ϔ��%�����
4d��K�<��ۏ�umH�>K�%�<���!�#_�K�|���i�<��N%��BX�甇��h~u% �����>Q))-*Z���-kJ����)hR[	1Lb��1��F��<��f�ľu��<JX|��������[��┄8K�_8��^|�%�]JR�P�_�J�K[����V��!�~ �!
B����6J��[JߔġJZ\��t�i�K������R�%���
q+CM|�'PZ��6����M� !�%��[k�j%�:��|���%Lu��SZ��������Ġ�IA�D ��(Z	jV�Е �!m�KRش�E1�~|��S��h[Zy�/���:��?8�k\BX�Ju�(�$�[�ĩF8�+m*yן<�|��,�y��>[n�א�)���P��)JSi[m��R�����:�f��ο6�T�T��⟘žI*I��B	R	j�_��~Kϝm��!���%�<�-���6��J�q�\K�BP�h|���&��\K�)�-�[�|u(K�JT��(RZД�Є%E-+B5)l!i[�����矘֒����y[8�5�1�<�'�S5+kZ�����m�ϒqkP5o���~C�!�hbӮ5Mi��:��K�����X�Ϙ��%�%���ǔű��iq-�-�����y�k��٘�1�d-'�m����J�B[bԔ��)kR�B�B�|�]Z_)���A�S���[��[B �8�����JJ�B�ZR��IBP�%j!iZ֓�k�m���hB[u�+q.��Hi�u-�!�T��1��yih�Z!�-�SM�Կ:�N-
J|��q��:�8�?8�HSk�i-5�k�)��Z٩i�m󏖵�	c�6��)�n%O�y���|�+? ��?<�kK��[BV�R����ulyS�CͶ�1�)�q��q�r0�P�R�Z	J֤� ��HZ�R�е�(B�J����е�(Z�JҤ�)JJ�(���T��IR��D!)Jҵ�Hjִ��QKBе�$��Y)B��kR��-E%jZ�BJ
Z�����%I)hJ��!ZД��Ф��~[mb�qD������)A�����Z��R���BR�-hR��	Z�е%[�!,)L|�� ��:���jP�ϝq	R�cϒ�Hk[C�%ג�KC�:mHb�q�X�ZCZS��XC|���!�>y,q/��_!-A��i|�g^Zԇ[u�T��4֜J_j����>u���HC���)R����,��H,�%R�!kK��	Z_8Դ�8��|C�l>Z�>J��ԡ�y�m)clS�T�!hq)C��u*|�!�G����6Z��kyġ�-!k)
BX���RV�%d%�QE<�)lB_?%-i.�����q� I�B�p�-~BV�A�5��C�ϞSjB��j���AO�ǐKMJ���Z����<֥!�-�^y.5o�y	B���HJ�Z��%IJԅ��HKf���Jb��!�ڗ��:�>[J4�^R��K�[B_:B[q�!�KjR!([�4������8�-��=�T��>[�P��KkJ��6�]S��CZR���%-ź��R�6�N))|��[�u��?6ũhS���1IBC�SjKm���c�:��6��M�����:��n��<��[�K�ǒ�1ǐ�qo-m��u�j[�8��Pǘ���C�-גS���ALx���\t۪m�)u�V��?:�򟚍BbЇ���yjb�uKA�ئԗ���~m�Rĥ�qi-��Y�,y*[�K��Hq���^R^m�a�C��f�S�ub�[kR)���u�	u��n��lq��S��Iq�^JP���1o6�ym�뭡km	c�K���]`�:���B�u�Kͺ�d:�X����miy���m��-n<���6��[�?<~u,C��b][:�%�6�lymM����?6��1O�~ZRƩ.5N<�?%)c�Z\b�~y��1KR�R[��Ko:�!O)N!*qM��jZ�JQ�p�ʸ���ۧP��Chq�ChJRZ�u*J�R֤�N��R����IqiBP�N��[��J�Bֶ�[\y��1�qLC�BB�q6򒕸[I�bZ�T�ugV��:�Ҵ:��n�!�K�p��bPbң�:�6��n���B�kk�ĺ��BM���C������RZ\Sm�۫bT�u*K�S�:���b]BR�S�<�y�-�C�6��%�:�lu�1M��1Sĺ��Bm-����n%Q/%�ug��\u��p�<��l�ZqM��:�\R��hmIC�V�֥�Î!�Yռ��1O6yĸ���ۊml)ԩ���uo!�J�uN���8��<�kB�yťM���:��:�έiq)R۩q�:��
u�R��[h)(J�ԭ��璝~[�<�%(m��~CV�_�ƶ���-ĩ����C�	l�4����ϔu��ϛx��R�-h-E�	Z���jYiA
Jև�%�b�!,|��.�K��P�o��/�?>K�A�8���N�I�>|�JTS�$ۭH[��\c��	Z�:Ԡ���%�>Z^Kh~|��)/%KS�u��K�n�Ÿ�P��A�kAo-�婵��hG�!I-	~B^J��%*B��S�Se!lSg6�!f߈I�6��u�!J1���Lm/�j�b�ӏ�$�_�%	Rҥ���
R�!hJ���F��1ka*RY�ΧLbO�5&�Z[~u.��1�5m�O��V�5��yZ�|��/k�%��䟐S��6R��@|�֗ϒ����%�����ߟ%M<���ֿ ����+�)�~%�_>?<Rb[-�k~S��R�j�u�V�yjCjcŸ�矔��(J~!E,��E��Ԃд%KZ��!D,�)%)R���Х))J�B�ZԔ!)KR�$�ք�BեiRHRT�%*$���RHJTBJZ���hBB
J�%HR	(�P��E�jQjQd�JJZ�!kB�RR�8�8��%HylJ����:u�&,y
)5�-Rc�T�5,JԢP�-�(R����%kj��)�B�Yls_��u	~|SZ~~N��.)O)ձ�?<��-+y�)�A��8�!	c�����	4�<�:��),u��]R\q'�KbZ%ԭ���J�� �)��B\Kן>q�B���KB	$�JBV���Ф(�����%,>CjK�的4������%� �>c����|�n)-�����bؗ�>J�)��ۨ6���8�α塋Z_�����JN����/��-(Cj~Q�!/%��ŜB��8��hA#�M1亴�!��kV��%��ϒ��Z���)��[BR��H֏��m��kKG�K��Ix���~KϐKZ����[Bpƿ>u)!+BR��J��QjZ���E-�V�1�B�c�R�Q�i-����HZ���%�Hm'�yL4���))|J�S��_�S�ı�8�ƺ�ژ�8�jq�ߝq�o-)S��!iujS~yKS���q��!D$RP���)�<���uǐ�h%-jS�C������ǐ����4yZ_>K�q�A(wV|��T�����Ж��^~I�6-gψA���!HRJ)jB��Z���m�RԖ)+c�丆��Ʃ���~|��S�K?%桨V��-�^y.�栠�|��)+~[��.!��jߒ��{P�鴾uK!�:�T�|�iC�K�-�S�~C�|�F�q�)�~J�b6�Ї][��~[��Zco-ǖ���r�yše��)B���ߝb���S�cQ�c�����M<�^u��t�%��~R�@�N���!O%��$��J^j�()JR�Bڴ�(Z�J��)H$��-	c�X�SS��u,լ�5lH���6x�)��!%��?>S�-����:�<���K�P�yGP�Ϙ������qS�ڦ�A�!�|�JT�1��O��m|��Jq��S�??<�ڳmy�|���u�?6�J�?)�bҕ)�~K�~SS���_�mh�����婫RR��hB�RJjR��-H-hBV�%*BT��I)JY
Z҅����%JJKZ�
)J��(I�MSRYR��)jZ���ZT�ք�*B�B�)HZT������[R��Y
ZKR�IIB����~Q*H��S�n�+qHB%	R�c�1-�S����.!(Z�JV�����hJT��()-�R�-(Kc_���������:��?:�J��������N:�����������~B�6��Xļ���4R4���1琥,�:�-F���)�|�6jLm*y���P�-�u��Hi�ҧϒ�?$�!���:��R����PIHJ��R�)��A�,�!l|�6��%�Hu$����C�J���.�^y����:�cn����)&�K��JK�)�BbS���o5	c�Q����_6�bR����))[aIq���S�F��K�/��P�խ|��P�j&�|���[~|�Ԥ���҄���u	|�5�k^y'�t�Ρ	c�R�\@�.%��Z�TZ��թ5��)hB�)h!
J���KR�إ�l!ic�����?("�y��y�%��X|��A-kR�!N�mj�ϛ|�<B[>B�J�<��ߞmo�6���ҷ͸�qļ�8��Ա)yלf�n�K�:��n����V��O(�����QIBҔ:�<���-��ƿ1/��<��q(Z���N�n-H|��k�S�<�%����y�A� ��u��!�#?>JJ^)K$�ڴ�IB������)ƭ*c��f�|���!(kVk��[c���bu��ZX��*םS�S�j�ז��!/-,m��c�a�An���8�-Jc����O��ߐ�B�|����%�_�A�SN!��K�RXǜA�1HR�t�_�u�6�����8A����IJ�Z�[�%�:�ߒ���c��Z�bR%�R_8�]y�甕-Ha���Zc�Z�:��|��ǔ��R�)JR!kZ�B
jP��jm����Z���%lK����%|�%ԾZ���Q��!��bX��1j��ϐ��������]BƠ[�)�jP��͡Ԭ�8�h"Z�~|�Ч�m�y/���)/:��9����+���k��z꜏p�M�������sqf�j�������|A3��ٳ�h����>k�>!���si���쌲��[
��F�M��l��}�k{j�Ž������iD�b�Vm�RkQ+�
��EKVFYIO�
GcQE�
o�H��5f!�jmcUSm��eQ�����a���ʦ�ҩ�lj)��Jl��k�Z!�ݶ4E���X�F�34�ic4��[3I��6j��jw��پ�7km���M��l�@wX7�%�$l��5`���X�)9��2�x/Z:�1�c��u��erX��ԭS���v1��G����M"Y��,Ć-0hL�ZY��Ì|�c[ƿ{��[m۟�:�����Ǎ���+��`��_�c��N��~w�t�_�"uM\/*a����e��п���cg��������d�V���[.�6]o!���?���69||��n���wޝ^�q���JP��#�澣��G��R�=�ie*�?&Wq�2��(��22dY�h�����'�e���?���=����K�&yt�G���;n��n��=g��t�o[�;k�e���w�U�������~�+׬�����7m���s�R�ݵ�1Y�7�4:,�&�����7��k�FF�I�����5Ŕ�'#��[������r;U�OQ�O�~��xbf]-z-��\F�qa���4Ռ�0�v)��c�}Z�N�c��;66��q�2!��&��M�B&D#BdɖȄЍ&D&��L�L�ݮ4Й2BhI�	2[!l�L�Bd�M2��2MI�B#D!L�M2!�LM	�&BL�&�LL��Y�Ѥ�B&$ȘD�2&"!&Kd��M�F����	2BLI���$�B&D$�4BL��M		��	2!4�L�dY�f��L�F�BLI�B&I��A�"m!#d�&�2&$$Ȱ�$$�		2&$$�d�$�LHĂ&I�&$&�&D�!$$Ć�6��3H%�F�	1&I�Ch�ilDbF�`if�6���Y�̖��̓	0�f�fKlifm�8pi��,�!,�X�,�L�d�m�Hn�1��!&$Ą��$�l���!!�ę!!#i3�v.0t�̐��b#m!&m�d�� �"h��b&&��"HH�&Ka!&$�L�LD�L�LH�A!!&M���1 �!4��5�!4��4B&M	2B&&��M4L�M	2BL��FM		�=�ppL�m5�&B4�!&M[&�2L�!��[&�!&M�L��4&L���L�L����14"4�M2Bm��2hD"	�&D"�6���B!l�4�Bi�����Ù��ɓ&��"&L�&Є&�ɐBi��&Bi��	�&L��Bm24&F��!L�#L�4Bd�[&Y�B6�&�ɑ�Bd�!L�L#Bm	��Bd#B5�4ɈL�d�m&�3Bm4�2d&L��2	��p�!	�M��5���2L��&BM�F�d&�!���	��ɓhBdh�hL�Bm2b!1f�Bbd!14&L�M�	��ɴ&�L�Al���ɡɐ��2�6�LM4hM�CB2i�e�m24&!3Bi�4!�6L�B	���І�4�!�Bh�И��f�	�2Є4��CL��kdmf��	�Bm4��ЛhA22�6�M����2І��	�d4#i���&A	�h�&hFL�i�m2&&M����&B2�&�FL��6�#hLBm2l�l�bd4!�F�M�&�#hCL�&�m2b&�LЌ�ɓhF�CL��Ba26�CL���	�d�B�@�	�dl��	�d�Af�F�&hLB2d�4ɐ����2m�1	��� �hCL��@�d��M��Й�2��M�d�21dɚ�&ɐІL�Bi�dFBf�2�ɱd&�hh�M����L�hF� ��L�l�4�2f�	�ЛBfL�hF�FBl��M���LИL� M��&i�&���2aɓ4&!L�!	�i�Bbdd#i�d&�C[h!6�	���@�4!2bd���0�6Bl��d#&CBl�0�d&ɓ4 �24�&�!�2�&�M�&Ђ����d�ɓi��ɲ���&��M���L��LL�	��4�dɲ�FBd�ɴ#L� �m2AL�	���Ђ4hM��!L�6�d�&B	��	��&&M-�L�L�hA	�&F�M�	�&F�Ѝ22i��f��2dЍ	�&��2i����6�M	��k��r\��YI��ie��t�M[Z[[���[��}���O����>�"��&��a6,��9_2y������=+�9�1��?8�K_��y���O9�	���\��������Ѫ�{���}�����~��K�5�S����IJm)��-e�z��#�^���=�l�����S�?qԻ��<�P�%�I��=��](�}Ն������o��FcЯ��5�kcƯ�r>�����LOA{����9`�<���S6.���޺��뺵����]��3���b�|g0��2�n��zS�ӖҥJh�Gª)O�|gކ%�/����Va�Yj�=�Âvrb��N%׃A�h��q#�͢��{K#�;T�,Cx���q�<�E��,O��)*��0�����ΫԜ˝F+I�ѕ��T��64bj�ib��5^���8�YF>*�j��-j�kU��{u<.tr��t�u�1�&����I)M�Ծ��>��V������E)����R�O�eV_,z��uR���-��9���?A���s/�y�З�^K�{��m-�b^��z�m��e�2�I��]S,�=������i���O⹧�OM�S�~g	�U�7��y`E��m�o�=a��SD}ۇ��K���O�_���g�>��ȼ�Σ�?Jt:���\�#��ȬX>A�Yӱ$�4�Gcn2�ǝ>u���`�}�0�����O��bf�n$���u����r�N0�H�6��oW2p�C��s�;yu=�]����}��h{h�Q������MG�69<XOAb�V�x�^��Na9����ц�s�;G3�82�)��+�|��fZ8�'#G�����H�y�>=�g�>f��>���^�K)T)���[r�}��}5������rL���ю���W���������j�G���3U=�W>��A�9����M�ǲ5hMӖ����Q|M�=W{���H�
�W 