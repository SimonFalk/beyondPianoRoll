BZh91AY&SY�i{���߀ryc����߰����a_ �}�P 	
JE@( � D

�� P        � (  ;�
QTzP�UBJP(P QB�E 9��  � x]��=����+�{��<tth�Av�N���*�@�O�����y� t������ l8\ �bv�]�U�#�   �T���ޖڅ�ޜ���#�mK�Qۭ��n�ޛ�L� T ���A{��p�]tz;�����m8/n�� �=ۘ�h8�� p
��w��:ӈ�{8������ܥݜ�^�K�=�!��) ���0[����zr�vq�m��u���=�����=o#8B�  Tp�<vz��ηN����^��m���i�{d<�\�x&�pT�@(M�6��6�o<E���Ӗu���7���1�����s�J��   XPGow�R-�����pհ�;��j��w��c��s����ݷu���`�gx6Nl=uM:���@                           �~ �&��6�@   d  ���%*���	�L  ��U)!M ��24�4F@i��jy�j�!4#!�����F� 4��z�Uڈ�&L44���
���@F�4hL���L�hM�<�Se>V>c�����ï���W~��66ٸ#M�cfٽm��1��M�m���m���;?�q��fm���N��[�o�{��v����q�x-Xݺf�lm����xt�ÇWct��f�k3��xh���4Y��7v���fcf��g���^��s�����~|��s��__���cl�-��������|ۣ�ǳ�x�W��Z�W�ȑ���?V��������)J�5E)�S���P������NZˑd\�2��I���m36)�p�&U�+A�;hZ)y��yd�a˹�B��)��%遷vs��]\���wQw'�b�mf�sm��x7��&�m^�2��mL��iז���4Z�lIv2�ù5곴� ̧n�ٮ�8��JT~ד�/q ��3\�n�:N���5zN�͸Զ&,�н��W�b�b�bx�ݨs��*V�H��8��*fj3yZ��[Xf�љ�=�ʳ)��Pr.(���)��D��xX�L�Zp�b�F�Y�c�7
� l"����ԻԌ:ha%+�oXȥ�Z�0�3j^jd�B�E�����n[���B:7A�$ǳM�F,UXK�d��9!�>�m^�#5�V��v&e�i�q��p���5T�3��)	��y�wU����Jo\4��P&��z-��sV�0\3k,�ǰ��$}oD��^��ݫ���.ȼ�]�y �)��L�z���[n����fn�V��Y�*��`h��Ŷ��[L�#J
p�hn�[�u��BD�g�.�%\7m��f^
	�ܳ*MY�{�22u�a��{��H2�WB�tԡ�fNKr�aB�OM6,�F�tU�,[Xt��+s,D�X��"�G����ۀ�otS���#[�2D9B��f˚B��͆S"��e�C2ae�IPƳ�be)�(A�22�[J������c���J� �¥��,�.h��f[�vr|�%�w,�5�"�R��$Px����Icd[B �V��qbe*1��4b��זR;+Crf�iXT�r��b�![PSU4���5��[��g	۴��\C3�Y�;�fE���vA�T���˴�ջ��k��j��r�jg/�JU���ʊ�\IFq��k�=�+�cPu��Hv3[�ѧ��԰V��H��E�&�����wq��īm�-�n���0imY,����M�b�g�UeZ���&T�(���`��pᠩ�tˍ&��7�M ��_�6��d��V�+�P#X����l'&L��B���D%�(M��*I,G�H'��\��q�c���h|��jԩ�-�Z�J�2�f�`,��4��˨.�J��`Lb髚�i��!8�
p�ƚ:����Xum����X�T�bF��ڔ��Fm���aY̲]V0��%V2C�4ꭷ�[�a?�H�:0�g03qA6 T!nc-+�)�ߌ�s���`݀\��	���k��
(���x�\��af�j���Rb{-���4����Ù�З6*AXD��T+m�P��WT�T�'p�����t3n�B��.h��g-�y;�b	��'�m��c77j�+�6�m��:n�*�jY�Ȧ�CYǢ�Y���� ��Q��F��iQ5���%�.]�2P"�`7�S��#��p�%"n!���l�h�ڕ��%��w�ݚ4��6����츛_n���5;�w^�M`�����\��8K�Vٴ	�p���x/w&���s\�E�W��%��d�����V�7�^ҹ��c+<�T�*�V&�h�r�&�-a�WR�Vr� ��{��o���B4�3w�f�8+3)��Ӵ5^�������u4�n���0�m]n��Qs�����AM!�q+$�K�8\�`E�<������Wh]�d��/.eE��p1�܊�n�d ��2��w��ͥ���Ŋ�۠5:՗��n
�*Ԡ�� ��l�Nl{+5Q[`��*�jjǯ�#�R��t���G��W�j�t�GWj��0��̒jw%�]M�Ô�9�l*7�j
�V�U,�rY�,��qnS@�9�MR�8�n�a7.�3s�כc6Y�u��+��T3(ݗ�l�Zm[�y)"V0�K&���V�и��p��EDe��*��%ֽ�*7Vv��ʶm��=w��b���S1Y��-���MxIA�K,�G!Q�)��[Ltm73f(��c*�ٴ�
h�*�S�:Z��A$���̴�5�&�Vb�Yf���+���L�r�@loe�y��|.Yn4͙R�-�W�<�X�(jݩ$�4*۠�U֐n��A�x���+�5+n}����!�9��4n��."m�Y+t���˭�}$�-B,n��@A<�[�2hР꜅�|��f��m0�Va�QTme��&����t��z"����2���ה�˫�;�/Xm���*�)])r8)ly
��(nh�oM+uV!�[i*��lZ���4w��rJۡ��gmk�F�)jipb�沌,�-�Z`\ř�WF��ZpM�akuV7uE�
������(�˷�ˆ���{�"�'*�A�#h�\-eԹZ�9&w�6��Na!e=L��[ԯ~6̭ Ŋ��]iZ��sD��.$Q�Ȓ��5`<F�/si��m7�I'r��mc��E6�KܖDlGr�Y�(��gK��]93�de��,D�L0;T�����fXj>z�)k���X�L��n� ��@�L©k��"ͻ�T����!�X��}7��Ř�)6�:�Z�+�&��x�$4�W8Qu(�A��um�f޴��䨲`��� ��)%:
�
��T���A�A��2i�p�y�,�P�pdV:�vʵ@1�Ay�9M`��&q�pg!!JnL]�TDӗX��@e�ee���F�'}+F.��[h�6��S+��Z���խm�0a���iG�+)[��pT�]�z��[�f�k�*� eVi�b�ȓr �]n�+3C����E*w-v����=��n�#�"�c@!V�� ��YnK���ӿ��G6���[�ALb��(�!)�VX��β
/&�U�u�+a˺a%]e��Y�mY@�wVhܥtZ���ʣn��ޣ�\�@��gpk�.!5�fA\�)E��-���K�B�7 �j$�R�naz�[��90�Oe�<V��4�A��L�T������/���$-�!�2h�Ź��޺�d�+d��6Q�7�]]�NVV���xuC�@�DS{Q�EKS�n�f�Q��df=�X�i4�K8Z�2��M͂`$�
��*�Ti�b����	��6M'}[Z��7����)�c�r�����g��?`�@#�����h�O�ۼ��n<^�ϛ��r��=�9y������Ϸv���������|Lf��5]������ю���Bn��a�n�=knۘ�y�ň5�w��u�m�n�mv�\�����t���q����axU�`[�1�Ʒ�Xoi���I�Շ���>��	dc�+ZU�s�p�k��;x.8pmї��cu��8�����Irvz�����['>mņM��T�+Q�`�"UPq���\]����?<�k��r�&�W�(�MI�.���f9 y��Q��NC�O۴�w��\<�"�ks��FC���X��񭵪�n�=���ʹ�u���l/m��lt���ㄷm���۶�kk��x�^�5f��S���s��^h��ƃo'ny�>�:�૏km�̮:0盟gc�������I�p�^�֏^uۖ�ε۱�d�`˳q)p]l�OJY��,�9�:@�ݠ�U��s�p��KɎ]��pv�{��[��=Vù�7������HnS�ƍ�A������An���;<��}��S�����m�燱r�7P�k�]v�U��؜ch�e{/n�����N0�A�Ys���p��!�ÌV�7��v��v�)�z�c�ۮ3��.����8ӫn��mC��ڣ�R�h��;�N��N���-��T9��۲<n�r{lL�.7c˰�-`E�	3�u/���L����i�u��:{m�*mfޓ�s7��Oe;8���P����z�n�{b��KعŢ�"h�^8o$i�J�k-�o]����`����kv𸹅騹�;��3k7r�+���%�����&V��ڼl���']����a���I�i}aL%u�أ!ݵǛ!;{��}���R��ݷY1˄�κ����ǌ���Žq �@���N����ۇ��PjwZR۫v����(m�n�;D��Nn]��Wn��[�}����$�b십��N{~���~N���>��.��L�v���o9����n���7㭎#�������ٺ�qգyM�8�u�i��u�,�t��E۝b`E�#a�]�T���Pٷ�m�z͖�pj��z�.�Y�^x��q����Decgy�@��6s�6��\;^c�˭��r�kҝ�{t;� l�Y BZ��J��=�􉭸�y�y�t�g�F�f͵w9��z�h��Q��&�,��mC�8�vᬙ6VY�jݕ-Ag\��7b�C�v�k�m�x�x;d�1v��v��<���;�u�ƪh%�88݅w�eÓ�<�������W�>��n۷�x��ȡ�u��A�H�:^�	����dz��緍��^�EJ����M�\}��r��D<�v�n�y_8�A�����e��Y��6ێ�ӗ�mr��6竫�;j���#���KVۃ��i�cal�����\�z���퓄h��t:DDNPT�R*�Pk+Q��ss��Ǥ�m�vڳ彍�p�[�z�v!��B7r�Mk�U���E�܅����n�{�-GbW�{v�F�ٓs�'n�*\��t^L��</n�vA�Ӽƛi�a����'@P^d�
�ݧvy^�]�EY.Eۂ��n���έ���;gQ���Ŗ.��;�H�ۏts����lk� �n��x����"e��7=�g�S7S�6�,[�\݋��Φzl��<�	��h�q��٨ۛL��ݰ[���:ͮ)Oct���\m���R^����Ӌ�
�8��v��8#��;�㭸�X�f�$dc� l��<�ƨ�f�#N*cm;V�筣{�]�y���ݲF(p8�x�/qݛ;��:����P��l�8¤�Î;�OW�-q�+\����U�ıcQ!��&�*͘7�����^S�ݗ%�h{fpS�ۣ\uk���gr�q�p�M�cN�o;=�ua���7�+�N����эz�8Mq�-�������X�|���\\���ڙ�玞��q�v�U�]<#�k͐�<�8{m�G�^�j��]�WOn�vlm2�l�ҙۧ��n���*i�-׷&p�8g�v��m�n��m��5�75
3�ԂA��A���/���=pv3�Chw�<L�b@�s�-�W�n-���r�����1a�NOk���Љ�_�v�Y�8|�����;Js��s���mC���[�ͳ�Q����=r'c;�iݺ5k�n�-��W��g��ڧ�amr5i�q��͞&�ݗpҭ�ۍq`��N�����&Su��۳v����5��p�c��b٬�Z7J\��e4�o�=���D����fٶn��nwM��q�`m�v������</?a��{�>�{�F�9�MΎ���_��O��߾�B?�s"E���U�e\���#n��be
cv4��Ϝt]C��Ι1��a�Y��4n�`�!7Kv����BdwQw[tzuZ��x��E�q�7t�0]�yX���!�Ϋ�0�
=z&����5�����u�ZK�^k���Fѡ���!��0%3&%�gT�h:�ϴ���q��k��� �g}u�hsl������>}��S�S1K1�{��d���i�i�<�o��i�ր�"�r"�e�B8R��qaL�Ra!��f�GE���Z�2� 7ӰҊn=�W�,^��*��T�HQ��'��Tc2�?ob������B��hS��S����\Ǖc��naκ�au�͑/j�j�;y�_<Vw2Y�Q��0m𕭅kp�וS�[���q8��#,]Y����맼)��r�����7&���Y����T%� -꽭�W]� ڜj��7�9�=�@�0=ܔы��=k;F}*of�#s�f��٤ET�ҙ�lu�s��������PI�s4�vh,��)j"��W�n�Z�D"�J�e6f}�I�(��n�kȌ�ne�=�[H�r�@ګ�3�s��R�3����e��#�ΦYz�oo;M\���I".\V���f152�ڡ�T�!��6V�p�S��Y@��y�dݣ���oN�K�0��������4��s8�C��f��V�Y'_P*��^�˦��Y����
�+a2�r�ebؑ5xC�hP^��)V'��
ϻ��)�����fV5a���Y� �<G&qm�k#�!�H�h7���f�;A
�4�XM�8%�U17t����R||)�K ��m�b)�e�T��6e�����m��YyZ"\�T�Y��\������wS���2�&6`"�k�@OYK���Y��Y�ʼ��t��j��l\�;s�_n@s�zl9Q��2���_^�Ko��¯Wːأ�/q� Y����u��.��Q5�1�Ʈ,�5���B���0q
x���YkK��'��Z��.�C��%پ[s���<8+��7�XjH��D�}�ZR��j�{�;4�G4���a�{���^��O�k���ޒmii�n���ɶ'u���������>�R�0�|���s���0�^X�y��ʴKͷ��`�f��83[�MU�R�8���Zy�����r5�B�74I*C��a�[�m���B�3���8щuc!�3L�<��P��Ŷ�*z�=gK#i���r�Mĸ��Ɲ��c
ŸV(�V�N]�6��i�ur��n���+�3f���9Y��i�·2:�t���̕�]��2�ڪ}����.:(c�S(�#�n�ɠֲ�wH�����
c��;�mLҝc�jkEԧh��H�{oa�t��c�<���ʤ�2�oa���I!��V�ctT���db}��[����ٷ��h�$��$����n�q��`�PH��;t��\>�ww����:��b��Y�-LP��P%�5W�[�ڸ�Ƽ��,XU�C�!��N�;�yUf
n� �nƢm̈́�F�Aٓ;�.�Ѻ������n+�;�tWyǍp-���,K�ܻJh�z\*ҙ��/q�����#+&+/1��
�0JΒ�|3�;;.�G�^�2�d���
�p�׏N�C�Wp�ǟX@�vk.����,+�'Q[��J=��}�+[����[2��T�;�0���z蜵Gn�
��+fFa5T/6�AI�H(i;R����p��**��Ř�SKk��N�nv��r���:�>����\��nN��%�+i-�-��PӘ��VT"*�3�H����+x��ս�6m\S����5W��C���F!
�1�)�Db��R����SQ��]�ե���A�q���s����,3���db�'�.�x����:kg�����М=��2h���o�u���Їv(��/��ł�ڝ�1�Ǌ��.��Y�MB�`�gG%�8N(u�Y��r��v���s08&����$�b �h�oF�wo5��1iIڱl}��u���f8F����DZ0��x��#TWu��.���(Mum<3���ƀ��(Q��|��Y��Cu>x+��e4w�+ˣ�.eN�!e���*J^H;D�I��U#��RU�'��*0��� ��3 b\N�Ri�,v�b��r_[j\��&�b�
Ь�W���qv<�;�<��jdt犒6�w����9'o{S�|^�f]���[��ÛK9�g1�.]G�մ��ua�W�E��y(��Z���9V���/f!\�Vj�6�MMn�Tu]egr����J[�O;�0�Ǥ�deK�m��yO��GY�2c����{�� B��;f�����* )N��:뱚�W�	B�[J�͊3�}��s�EW�]#�u��V[f��'� ��r��^ò��b�7��b�+7n{�cM��ޗ*�����8_z��cr��9Y�n�bNֲ��G�г��k��L��;�����c&�Ӯ�$l�vZYEy'6�����=7��g�%���tY꘹�|X�ָ*�u�����F�rѷz;��]��F�p��qn��4�^\��-g*ۻY�%���w����ɷ�#E�Z�rk�]���lV�,R{�(l<��_fsF�"�Z���))M�^^P ��>{����7-=�	�@��%��1�	�wvy��{�sy�ƳG�*���6���Ɠ��!nT��Y�q�=���+��I��[��t���]�J��I\r�9UC)0u����l��"��G���Q�Ѧo-Sn�y��8�
M���>E��V�Ӑ^m��N;%f����3Fe��oeu-���d�p�ژ:ӆ�����r�fY�|l���c.����K���`r+-\������+"`C�6QeFm�8.V���gL}v�}S����=�og}���Y������!!'k
l0HE7b��Օ��"e.�w�a���c7%%(
�ײ4���W�����|sy�w��7#�up����6^N.�l��`������%[Ү���[��(��YX/FPW*����:�VW77A.2C��V�YX�[xkz��R�u!�D4s�ks@��mn�v�N�緱ӻ�����z��f�٬[Y�W���k�}�6����x6wa��z\����ߗ������̞���i���\��)�C�Z�m�
��a��˸b��x���XgP�d��r�@�v��9�\&��I����[�Q*u�NM��Θ6����I�tNܗ/FI�ƞ��<�v�n���]q��#s���9�Pv9�m���c`�7<��y�gAf����������x��硝t;;���>�u?Qk:�u�v��{!>/Oiìm�mԼT��u9�7���H��۝l�/K��v�6�]���Z��;��`��x��ś=s�a��eq;��������:8ݻ��׌\F]��%�`;Y�\����2����Mɻ��h�v�F�ě�۷gv�3Þ���u���)̶-�#���9��qu���iyØ;�/L���C��R�b���jr��&1Z�B�7n{��Od�F��^�ㆭ��-���i��2�[F�e-�.�΄-�q�rfkM�I;Z�P�(TޮO��\g��Ҧ~�4�$m�P�ak��ڙӯ7UZw�Ȅ��y��=3�Y��Λ�C6�}��n�-*$���>ə�c�v�!D����N��Yxq�-ti�V�1�z��V6�h��އ�b�^<$	F-�+Ss;�W!���[u�oi���7��׈c7���K��V���1�\���e+�׼'HvX���ӧv�|���[��6�Lu�8	ѧB��ج��;��T�uI�{@�&Tɖ���z�䲷#G�j�$$B�r�VBi�˫�R��!Ř�S�$�7~ֳ�w��kx���5��� [#(U���!�O-��n ݭ�l�Օ&v�9���o)�.Ż���XDo=�]�3n9Ok��nƁ��mj�=+FA�mv�K5ftnӎ�&��dUU195�T*�&Z�۽nG����&7���;r��&��=i^���_�[�_��%
��jB�M�7v[�>U5�J�JB�p�Vβbhr�*g�:T�8)�RQ�}ܤ��#�1�d���şD��ֆ��]|R�����e�%X��c�=�b�����j>�LWX!x%>��)[�ɸ�-����c-WI[{t�G�������C�U ���
@��x���ՎE{��[�7j]l� �$���74l?�t�Pr�~�}�Êq��9�O����t�f���_"*_r�G�*-WB)�n�aKzkK`���},@��+�dW�e�Cj�,8�Sʢ����}ԑ�g]���a�ݡ� Q�5HOBKt��*�����!K������i�=KS��u�,u�[�p��=��hL��+!�:&��Y5��o��v�
T� ��~�WK�D}��nCQz��yQ`V�sb������VA�H���z��;�鬻�s�O��Zo�qo�X�%�X�5�M�����]��\~~���&���I\��ս�00�Hz��_9]�/�h�z�Nu�� ��mp��D9B��S1u3����o�B�
Y����Ҳ�8��BW"�8H�.��j���PH������|zr�
A�*�b#�+"�¹.��Yı��)s>��k�f㵅6x��v0��c�7���[�e�C�T��u���Dbޓ�8�$�m:�<�8P�c"!��g>�ܾ�Tb�S���͉����c�?u���\)'���m9�Z��諵n����v�U&N�l�:�@�cgv�EŢ.�6�^�ێ���s�i�N�!����$;*?���wʟ
���ݗV�S�c/�+�k;���W�,��bQ��A���αg����]jh㉎Ȩ�]V*5\t�N}*�&bC������9���1���M�+!��C@ ���Vғ����	�� �����s�֘ED���Ŗ�U}� ^���CFy`#�9S��Ӹm�h>{A7���]�-�ѝ�ﯾ��p��jj �@�*��
�k��z�30�;!e�gh&%��jtP�#J�>`C�r�$4��w��Ф���H��nZ~�r�WNkt���U�����d�P�8C�B� �(�vڈa+֪��V�I�h$�7=������Y
�&��&+� ������S�Kq�=��ܥ�("����f/�P����z�K}Hn��`?VaM�#ڢ������0\D���9?|���m���:܋�0��!ƔI���ሣq|�*-��52�0��y�ɻ=	O G۩��$������X�q�uqE'
�qﺅ����Y�F+���,c����w��qV ��7J )Vf���6��X T��NM�`R��L.o��R�}�����B@��$.S�_ԉ	ӽt(8�v-M[aЋH��SЇ�2:hU�M�x�_�G7(�w���-����`Uz�/���]q��Md��,��J��+��.ﺙ��ݸ�ls�q�v���@���v�W�k�i�-D)�]�#�V*!�3��˥��"Ӷ��@K%I��|�&h|@�"�r�d���(���6��P�PD�)�"7s��G ȾӋ��|��3���O�F���4~߻�.M�#�ʰx�{v�W�Ew�7j�����b�=�nw����N���玺{B��I� ;z�d�jv�{p�=R��x6��헗8�m�����[%G�U_	R�hB�W�O[��Md�T涣�BcjR�85�VK���V����}#���߹��Fx ��1!g��h�{@`	"9Y�_b�w�5G9�) �:P�O$���������
��	��Y�j���\��Z92�tO�E>��L�R,%��ʊ+1�إ���]ܹs����HwV�8Q͜f#�x�u��GK�C{��u|�bT�]A`�$��ϡ�B��3s,o�g�.�ji�'�B�aҏ�O����g�fkM�'����K��B56�T�*��Pr�p�,o[ ? �ԯ��>�����v��:d���ي���B�0Sjo��Ζ�!�r�(h���ֲ�SmK�`0N_B�D��l�/��>������uE���F=Y��#�8nF[�mI��r�.�sh�;ْm�7�5���L���N����b���-�t��c��e٘�Ŵ��/'	�'����z\9��t���l^���c�*�7
=�3Ǩe�.�����Yl����L�<JŲ��0�+�T��+?)I�k48�H=��5����QQ"myyS�x�}]�x��v����u�^���,g-I��=�7#����!W���K*�:lR{����/]�1(ٚq��=C[��J&�K[�Ix�ۋ)�V@�Ԭ����}v�K�&c5\��¢뫳�����������n�{������Z�H�z3kk���=�~��ߟ?8CP���>I�H5E	��g�Ss$6ˑgh�)��=���ז�Xo��"㜒1n�Gµ���Sx;z,��V/� ��d�Wl�[��RGv!�<�V��Ekh���jE�@Vf��iI<9��#y}}I�t�J�6��j�F��H�M�X.F��jT�ĥ���݃eۍ�q�îwa �|:���l�`g���E�	f�	��	��Q˘ڟI"�z�U��9����� �wH݌�1H�;P���͢�-�Q>�����=۬e;Β�e�X�nQTtl�K*�V�f�j��{���(�ː�}��@J����?|>2���h7f���e�J�~���ѳ.�l�|{O��guEAI.��
U4�P�U�Or5wf���K�ESI/ǝ%P�[뤠�/��J	p�Ri��䤨���KkZT�*��U�֊�*^VER��T���U1wN�P��YS��(�Yi��Ruu�<Wkow���z��n�ЕwA%
IoW*�K�
�o��WT�%Vڤ��^s�s��Jۭ�xq�ru�圅c��m�ͺ����ך�.$��ֲ�V��JJ�W��B����1�I�R�5J	R��*����եQ���.��@I/cIA$��T�I���\���Wt��?ѩ��K՗#�"�i���_�CBL�@���C3�.͏�~X����U��RDH����'V�F.n�o]{�%�oM`�V%]�s��TPIW<�	R*��U�5J������ٌa	g�c�����)U�
:�UX�-�c;ZfVԳx���'}�Ŏ��0���vm��+��j�RY���[z��EI���m&�T�Uo�%
T�(%�����U�pd����}>�.�J�ҭ���*b������:�J��ET�^�*PT�k��-i�V%��T��(*��H� U�	TU:u[)(%
U��yu]�R-��T�xD�z(��t�K��TR��J
��>�����W!-�Q�Wp���_q�ڸ^_���i�D�`;�����*8W�l�b�e�h�g<��r���=5��5۫�/Xt��v�y�������n�0:4PM��Td,M�+�Q���El ��gݛ��O��jB�����X�i�����ڤn@իFZ� �8�E�C��:�x��qK*HGe��K���Rb_*��%�� �S涕�h*���*�o�<s��\iV�U�u��KU)��֒�*Y�$��m'T��E��^�۪
��:�ET��R�ZOI=�U
�ߚ�
U��;-��UKu�R򦘨T��*H).��J	-7I��MSU�5P�K�1���4��jU$�t��^K蔥�5J��҅U/�"��uk9�Q���n�=��Z�F�h
9��wڧ7-�]&�Uo�$�*�k�*�*_dQ���{M$�+),�쏰�Cj�������w�ԅ>���(X3<v��H�7�+�|![�{\�yg¨m,_~4H۫y�������os5ﶂ���d�T
��J�U��YN�@J�{v��N�%KU^ڪ�PQ �����R�:PI#�&mqi)5)WU|HP�)e��Km��Ux�XIZ�(��ȕ K��0G���[K�Ҩ*_%�J�[�����J�W�5U�V���Z��v��۰wd���G�Ki�~z�x;�G��uIq��yU�UAIo�R�*��tCŤ���Ix������	$	sΩA%��AJ��T���ZT�w��V�jH�U ��֕AR�ڨw�����U����.m��'�Z�9�]g�s��h�L�jr:��La�1�����#�#H�.~���3��t�����;r���t�
�**�i ����A%X𔫐Q%(��+¥�*9�cs�SN�Ē�:�U�����UAK�
���KDK��}���xPPn/�
%#��E����6M�i'f4ҥ�E$W�UPIk澫T�U��T+>�ȭ��Y��j�*m�[mPUVi�I{�J�SQ^&/�������l�_u��UW�P����ZV�gdJ�W��%
��.+4�i JuHR*��u
����*@��Ҩ.vl�\�;Lsfq�5K��k.~�$��}{Z{�����dz1f-�C-#�u8̹P
�֪�K{�{�n
j�%K�IJ�{K�uJ���U>u
Tmc��ρݰُ�F��"o9��c��f��(��$Ĺ�UA%�4�)U�\J�'AJ��"��k9�y-�]�[X�yYD�) UZ�U���$
��.U�H*�ny��hm%�R�:�UoR.����H,�UPTm褙IgM�Kz�:�Ir�M%��UP%�4�
���P��h�!��($����5RjR�]*�R�+UbR%����iB���P./�y���[������ݫ��'ae�� A����(r���%��q�=���K�lCh��8a*;j��GcCp����83��k���VAwZ�&�v��=��O����x��c�Ѹ�v�-ہ�!14f!�mR�U�Q	~8�(~N�3z2��6oz˺]�̰��IT���1K(2���"�U�L�,-5��b�X��J��J�V*Yˊ�
JT�i%����Bɥq�%�uUr*�W\"��t�K^i.R,
����xC�n�*�����]R�E� Im�H*��҅Uf��j�@f�����Ҩ$��J
��U�:N��"I��3��=t�ī�ׄ��B���5PI/�$�_ΩAWv��$3e�9#��rA�NE�I�����>�wW1���H�Y��I]3�e%��D���Ck�?��0���\�e��G�� �A���#�4�m�U7��7">�xt��Vh]U��EB��]�@쉁>Nn�/ 	�x������@ۥ
J�u�:iW�8��[ջq$�/���U-7H:�Wm+U[�PJ��Q*��X��U�*�R��:P���Yn�=H�]�I�}��AW��k�,SI11.�.c�+I�\�QU�:�Z��6���1�Q�Z�W,qڀ���[W;ҝ�kp���u��U�^]*b^�T���k�4����PJ���cR�Wz"c�b�앬�{Rr�h^{��7�����ʯ��bW�~�3>/]��ab�~� 	���n��z���E 2�+v��jyGx�NZW��Q�'{/>�4���0Ȝzڴd���Β��}�N�BMm�:l��/J���G���Z�k�־j[K�s�x_�4��Z=f3]/O\�ܢIEr^����2$���/{���[��ţ�%������Aߝw^u7@,���,�W,���Qu4��Pך�����{�\�v���)����ӭ��.�vQ��4U���x�z����l�4-I�8ö����\�Q�ɵ-��SSʵ����Ѷ��+�kX���ˆ��ڐ�x�bk����9#�Q@q��x�)MF!�ʣ�R��8 sd��瓚�y<�IZ�$����"��3���N�{�0b���G�R�=i�ʰ�[NiuT%(c��`�7I�|�]k�ঝQў� �.�}�l\(V�ti���qz���F��ˏ7r�Ϗkw��&VS�32z�{Z��|�_pK��̮����'��YmKt���]�g
��t2����p�q'�w�ا�a�	j����e���Y}`c	a�ݍx�q���k;bD��vs�W���-c)����Zǵf�̶�i�ĆL�{�.����K�s�a^�h�q�%�j�(`]�YN�N�����Z�a��S�¹f��2��뾡^�G�8\B�gwz���s"�~��#�\��x?vm켭���{��cɹ#�����GTl�_D7vkr/Z\snEn�
�������d�ȋ��M�8�%���U�y��k���vTK�S�]e;7r��;���w�S����%�JYc��
���ܙ޶|!c<m����'	��3[mn���'�+r[�:�����wC�]��v�۹Qwh�le�\h�d!%�s�sc�����m��Y:_<��g��`݃���k��v-u�ǈ����"�s��؁�t�nm�r��g�UN�*�ٺe/9�ٳ;n��vE{��%����曧���"�$Mفۚu��#Ǖ�����nn8^ݸ�9d�}�>����v6�si�v�msE����s�t�	����!sӗ�j簴�1�-��nI���y�T�������Q{{zl{`<e�m��S�;V��kؽ�;�:G���	7vh�v8�Jv�&�)k�d������Kn2��f������{��s��t���h8ճ�|���T���6z�y���7�ۗ�*<n�B��
{[t�m�<3qM���m����!�p?>�o�s�ۏ�k�'m�9G�]Y��ͬ�(cŅ�|�4Sp^��r�K���T.1�-�ѡ0���V�uf�3�s�Gh��	K��{�XNZ�^QÅ���c�U\�m��'�y����ju����8�\��w�Y��l�KF�!�wi�[C��찈׃�<L���l0���w V��j�v�8��)i� �r��N�-���q-�S;@ʺ��%�.���Z��Y$���`jRm��{B�&(���HE���������0����ع�Q�e��rG+���+�
��י���y��gp*�3u1%���IQ��k�ګ)[��ԍNH�R.��L0rY$��(��W�˻`dƹ�cd��nuó�6�ӯGI�7����|�;����켙���$��,���d����-�v���	���č�VY1m�Ug�w9��H�2�^���GG���rVG���Eiu��o�j
��j�q��a *���msa��N����ZJ�|�{��������� 3)�=,50����VS[�C�8��Ug�݂w��,�"�p�]�ga�[X�N�>������Ro���
i�{�3)=�t�gF���, ]�ڂv�ղmg.�!�\�{��;�^rި>�I=��~�W���5^�Z���4�����ӵxQ���ygm*|���!���o�<�*.�T� �:�N��?!��H����|#5��vh��bڴ;T���Q	w&}�rY��y����ǝ�#�:��i	4꽍��+I��{�$y�k����er��M�&�����IU��ۇ���[����~�|��Mg3]��OzxBy��.yפ���i�Ks�4z�K�C�����,	�F��Ӭ�+�+}�_a7�{�g�`If�����բ�靼1M�u<� 1غ�ӻ��Kx�6v׾h��W����\�Ʒ�XL�����g�ޮ���|���V�N�4902\B��b�EP;��s33d!�>x.���0���\C3�p9A�7岄հ�y�z��$��,J�}��V|H'�����1��`O�=p/�=�er�՜����H�q���!%d���1���F�.�����n��.�2�x�Gw�(3��V�M	
0
�^R�g�!-*=i��{�fEd�3N����u	��'+K�;t�t�(�,w�m���dT��Kd�ˀ�� ��գ�9�����.���Cy%��[A�ˤ�ރ�p�]@����k޵f���2�o~Bb3��o�ݹBѼ��v�?8H�y�}X��^n��>��.�J��6t�S�zzj�u��!\���ǠaK�)�x�0��=�g������n�tlS���[.�6\u͖��c�N��#�M�<l�ٚ��m��2��VM��n��r�n����Z�u��� � W���O�SNl���v��M2؝�?-_K!�x5Ǹ���R��TQ��:�c�9&��ۗ$-3�ރ9�_�Կ]���3v;CZ9��V�k�ϛ�n�_#Y��b&��L�g�z*��;3�Hu@���q�Ms���h�C`�)�e�"���?
��U����^7S���M�1L�V�["B�W����p��y���W��^tN�ȴ�{w���ٛ����$����}B_�\�Z�5��8?("'b-BwLX�`�iadԉ����&/�9-�����.#z�uyB��{���y��	n���W���T��u��D��j�:�h�� ��G��6���7��	�s��A������
(��C���sk�ۭB�1ZR�`�:љ^^c��닚x[I:־흄�"s<ߩ��.�p>0��SU�9�]��fE<���4���.��Y"͟O�G�d㺀�2xxA�n,��-���}'9���L56S�Qf�[�W����qM�<,���2�x��y�9I�~�P�8�ʷjog2c(�{@��1�c��x�����ݻp�8�^�z�5�~{[�a���	3������%U�o��Q��Y��=��E�w��+�h�H^�G�}���3�<2!1+APW-��;�6���>����=��c�?}$(A`�M>W�jଢ଼���G��i׆-�E���Q��v�h��Ym%�Ss\߆�. �x��0Ȅ���Z�.`��!�%�:���o���ﯹ����{�t��6��g�UN�g�ު�D)���oV�����k/ȕT{�ŷ� :�\Y�R��8P'>���8��>n����n�o�CL��cg��0M��i�u&�ѵ��ۓy�"�ڽ��|#{6 G�����������K��U*���[��֞�}I�y�cX�V\vnh��w=$��t��ӯ�^�u�7;t�س\�[f��}�����EQ�j�*�v��3ok�cx�� �G�̵��r	��y���lvt��ޣ�˄kiӼ��@������z�^~a����A���ri٣L�s�B����2(k��E���\rk!�U_74��� �/ɢ���X�vo}�uX���|��I�B�n��>�K֞e�}N�fǚ���[d�Ȑ�1&.,LDQ\9B� ��hҊ��0ꏵ���O���RY�v%?8Hϱ���zFڮ.J�zY���ֈ��(������mT�N�^HI9d�ܲ�"hd���[E``J�m�˩�P%C�n �TG��wM���%U�l�â���t��Q,��R<s�l���C��q�o�`OY�l;�M��s2!��|�ک���e0W+�Ē�[��g9�Җ!P���ѯOǤ���X]�I��l��Dk��x�5�㘎�@�.���0S�səPW��7�UƿPRY�Yg\�׻��JόF�C�ɼ��y�ꮍߒH�ّ!%�3��H��f����ҳ��̪�����`���.on��� .��	��Av��w=^eI��,u�cpR1����z�]�Ȼ�e���-��e�)V7�rqz7km�ª�V>��d�݌��3�iX눠����R��������Ф_yǐ���lb����ձl\(<�;��r���Q��hŘ���8K�$��ͫ�3�2k��/��]a�>��Wc{:U���Zr���(1G�@�q�屇X��E./'A%�PVp\:{�T��,_�͈�{����3�8̚��x�;Ѱ���^�472�]�3S{3��AN!���/�Ї�7�Ep�ߗ3>Qvj���
B2�ډ6����w62g\%SscRr[���T��ѭݘ�Բ������XU7�ۼl�X}�w�WLV&�;�ܟ=��]��r���j��
�y8&+�'e��r�H�)�$]�z�_8���s�@���tF�nfu��H��/F'j͐'qJҙa3���/teY:c,䱸J�P[��a�n�]���PǙ��]�\n�]���pbcj�j `�4���A�j�ڜ���Ԁ�.�+Ls���d��dEu9}�V�Z2��ҦP[ �g:Yf�a#m�\�f=젮�7S4셓��mU���k	8���
��UVe	v�rsK��[}�3]B�g�UC�<��~��Y�N�f�˹a�䞪����N/����p�U�G#�	"���*�d�&�2�'5�l��ɚ�S$�Yۇ�}楲�^�v��x�w!���x׻�S�"D�F���[���y	7͘�G&�BJp��'츂})��y��X�F��0�ˤ�Zᣟ��Ǯ��X.��Q�D��jR�CNPۀ��ɘ�0J���=�*Fa�������~�Z�Z�=x>�n7ݽ��5Q�b��V"���u����]؅�Ǆ/>�h�>�({�ʎy��� ��ߩ�ˎ3���#?8Hϵ��'i���I��Α�&��O<���N3C��#i�e��BLN��G
����ܶ{3��ǖf�+A�G�"q<�ڱB�o;}��Kh��-A�8ԗt�-*qȣHA���+d� ���+��]&��e��9��:�{r4	Ԅ��vz�������[��c�Ŷ۹�l������C8����s��;f7Von��3D�Q����й��7�e\R[⎲��ڜx���&s�L�Q���樎�/�:�z�5����3���Yi�`��j�L1����:��zD����O��l��E0,s]N�-@����u����g":
UF��}��qG����1��tm��t�s��h6�ofN8�~�BB�*	�cul3>z0�����=��Up��C�?A��U}��W�gGS9��ak�6D���Zh�c�����Ml�:���yt?"Id**��,��F�nQ�����;��L2`�����	=o��	����f+ ���z_[g�Q��i�ȵ�C�!eC��wD1�g��ԛ��{�$�6P�͸fEC�fw��)�Q�Z�f�nk+�~w��1f���j��^�Ϩ83�F{Y^�Ȼ���<ܟ}���3��DTs�Ԗ�L����)g���-�Lq�(��2s�9�?92�r"�J���N��S��΅)���{1x���k���#?8HϾ����tC�["LeD@��H�o/ݤ5�h��t�|��5�e]!N!/�[����\k]��2�6;߃|��I�;��������ٹ��ZCa�-]Є ors2՟ryP�>��aJg�d9�k����y�yR�Z�&X��v�7澥��O��"ߧ��P�w�c����۞��ң���n�i&�j�EIjrp�������	s]S�}��~$:[�`0�4w衔��߉���E���F��V��P���q9���:���ƍ)5���m��V:��Bl�C��_���gk�Z�^�P�H_�L�j��i�*��oU��i��E��Ild����^��σk��L���>r��R(�~A��w������
3vA�$�2g�8��KA���w�ߡ�s�\�����B��n�_l���p}�`x�M��-��Km���v@�կ7Z@����j��=d2!��n���f���V�@��0���䤮ϒ��gm���F��=��\R�k��j��e��B.n��=Z��'=����Ò��m70�Y&{��A���a�E7����7�1Ϙ�A�Hk$�����T��}�l4�I�0̡�[B �EF�׳�Ĺ7�ⓁB~˾}��܅�F�>���5���
$�E[םܺ�o^�n0�B��*�Ɲ���gM�Y�-�׸\�>����w�'����~z��z!��OLD�aC� �j��𨏣q��M�$|�R+�������ILgH(5v�Z��И���4kX���x��	�ĿF�?St,����]�G�U��"Ak�z�y���)L�k�����͆��&��)u�xC�	�kty�b�6����7�H�*;d����q[��%�HM�I!��y�z���'5�}���)U�}"q�Sgy��}p8DG�'�ٛON<��Hi�uܚ�3��x�3��B�-(� ��?Y�=�t�b�*qL���晢$�C�Y�S��B(ȱZ���7u*U��I�r�ߎ��,{�JA����
@+e5}~�ሄ��~l��Mß��IV����Օ�*"�ц�A�i�G�պ��0�+O�M�~��"�ߤ3|�;wq�[ɯRu�rF�-COt(P�og�Q�|��O`���5��\9#���(@�"��yrm|k�!bE@���br F��
���.�a�1t���M9�z����Bò�H�=�0���Ms�RFս����E��
��	֙ʵ��C.�޸�4��}c��V[YܒI�&�]ĥR<1��Z��x�&^Vqj�>�<�����k��,-5�t>��t!9���st� 9�җ$oV�=0rډ�#���� �/�TB�N�s ��1������Sa�Ge�3�7�$.����2����U�7�}��.��1��ǕWm�(�4]��)�db�(U�P�v�γ�q$Be˝��M\ؙ���Zڇ�c���e�h��M��Y*6L 2��'B�n콋�v�\�j)�\sog��{Ou�]ҹ��{q�%7 �$=̛cD�^TךͪWnÝ��Xë9�����]O���^_9]A�:�5s�y`lt���.{��R^�9w��鴏"J��T��v���D������KA:�hSi?1��t�ܲ�́�wD[sB�4C�N>�#X���C�R�]�,oN�v�;Ij�a���%#��iN0Q���u�c�i��$��͵yrVsU���.;�6\NL�5�D`�7R��4��C(�b	"�RDnDi��W��&�q�x�9ͺ#��mm0�U\
��mJ�(*�!L9��A۷fJn�$����C͙���t;��;oo=t�]��f�ǰ���I5u�ȾG'Hv�׬naʴ�mq��+�lEѻf:-W(�s��ks�p��]�n��ZT���Y���L��l,tQ�+�0�S��kg���������;v�U۳�uǧ��g��|ݹ6A�-I����/s{d�b��k�=��9�ۮ]�I�l�Z��fT4�v�n��rJ�U���]������;'�wOvN��랫�Y�^96{e�klu��ۏ'�4\��ՠ#�-�뫍e�����y1���I���Z�v��"���v+vS�i���:}[9��/+�Gm�8-��U�	��l�Ov�8�j�p���:^C\o �����y�=��5HR��/c&��|�o�R��˫{y�zS�ܭ�!\k����遮t�����N+9 �c.�V�ޮz=�y�m˩�V�f�S�j�A&
�nJ��|kUm�7i�}R���@L����z7�>L�to�"��C� �'6����*Y�M�b�BCSwy)-�f�;lvU�EU��sa��`Z��T�24�v����9�y���:������/U]�+�����) !��ACWw�%/*�Ǡֺ;kt�ɪ��]�--d�����#�g�K���h�ҳ�,�G^!1��QA��4737U�%F�5�y�_f�p\�.�w�_ ���+;1���ɶzx���m6�wi��w�s-��65�{T���s�q�g�n�dl���q=S����ss�z�w5ǔ�c�rg��Ǝ�K�\�;kt�_	0�l�'�����\İ��-�ʞ��W��t������Oc7�b���W�?"5>�����]��1U��M"\�)w��C�[��V%����I����9�}��K�n#�h/Sx�T`����;�%��IUs���(�|�~֪�յk�Q6{����Y'Sb�d���yKh��*)��+f���g�����76��ES�P��喹nռB��حn,���q��D'i3�q���Qţ���k�N��.I1��K�d2�y-�.�c�j�g��gx���R���bB�D�U�	Wt=]|�gM.�s�t�GP���K� ��%-�0����'�{.H�w�sz���4�M{��Y�����&�}>Vr�1�p^�?���q�\I���H[��Ez�;I����r;N2�YWq����� "h���q�l�I��y>I���H�Eo��Yg=
7����r��N_���q�<ޫ��8�?.�Q����kNB��Qܭ�?��m9�O�۳�K>^�a�e)=�xj]�Z%2̳t�X�f�ee.p�W�a�Ϛӟ>=;�)}@��I��MA�d�-���u���|A��&F����D:t/U�P"�n[�v}����C����F`��pj������k%�3�j����ZK/
e��G��]�n��fc�U�9!��^��l({Qg��6fE5� S�]���k�C�#���盫o�[�݈�F<�Î�{b� 
4�"��?
.�.���O]d˶��0c�_�x�fٕ#�'	�T��UO�w	���Rt�B�6����y�;������E$NG֤Œ�)lbGD�wkv�kXe&����=?D�D~����Ω�e�֌��i֊D1��z"��$��{)�ױ��$Oވ}�<�W�����5�xNք�A @A�+��T���E�G�O��39w��;�vW�O�o>��.�Wi�'_W7+:�Gܫi�%uö���X��ɝ�w��9C�[g���=Aƒ�5	���у;���񅚍ۤ��z�L���-�g��f92y�<K���]��}�\�R؟Dכ��Y�� ����;'+��cz���93U��78�L<�ax��ƞnݬv#����6K[-^�8;���X��L�H��|�#To�� D�~5�כ:��b����B��m�Wi:Qc���w9��	�u+"�	̖s�@��@���/��"jM���|��b|�mDCᜬ_4)��pl�24H2�2L8�dĩa�H�x�ɇkܯ�'��٪{�!8����}L6��'�}��ُf�^l-5K�{v����@O��a�|N�b�E�����L�3r�����/>���@�6uYdǸ��������&fނ|I�0�[�����s]Bt2(\�Hh�pͬ���߂ϰ(�8�>�#��Ɨ}�|~܂���ݫ8x�F��Y�-B\5�k=!͸k��E�A�I�u|43U{�?��V��sfXҎ��3`����b�%}�5�d���/�)+��+�QaK�5��M<~i�W��3T�����]����٧.�^M�܎��/�;�FC��n-�Y�y
�R+ħK�>�C1�RCE~���wq�[�v�Xށ��b��3�x��Rʪ`�^�/��t:��w�x���G߆c��!y��� o�<���$��Ⱦ�U��m<ԇ��*��.@�=O�;��Б'ԙ�Ś���k�*��B�cf�3>n���xϯ�3�x��H򋏏 $�u�)]�LT�ay
�ݝ�+!Hjg��
��*���ӷtb_�-��i�!�Z���8��k�!�)�X��z8�	*��XUer�89c��'v��Ymi��l�7�(ĐMkf=����1pl��%S9��}8��kH9���۹��uM��b$��g'f�Xq�>��jNS�ѯ9���y�r�c�!|*�o��<�V���P�$\_�>������ �	/o�0�+�`>2�'����.�b�;�gMˉ��n��q١p����Gu��ή��۫u�f1�)l����n{x½c[�7[��ۙ�l
l.��������e��^.�h��j^�7�FR^����<��#+dk���N��m.�Z( ,`��~f��5,t������i�|ǝ>�ˌ�ryP�#�p�H{|J+@����+��Ho�y
�E��I���˴��WD�e�s�k$�M1 ��4�H�l��r���3���f��F� �[�TR�LWh�
X���4����n��ω:�m��}�Q�qY���|�f�.�2V/[��lv��쯪��B�Z$'�'�Nk��N%�{�{Y7���l9-s�:M@���_yQ �}!z�޹1��(ϡ�X���g�@��F��ԇ�忙������$0��^�Y"�kn��=�P�L��Y�䞡�V��������.���2x4%�\S�.󠀺y������]DBiMo�;�L2 L	[1��L��'���� $�������x8��4-,*�� ��co��+j2v��~�^��.i�"�#k6�Z1.�շ�M����[i�}vw7z�ͳǮ[O�\I�'���<�/65=*�5����^��l��A�:m֬yي��ިĺThо'�42���vT��+V:>�-/�m��%�ݮ>�V���&�wL*-��S��-,�38�W�PJ�Vt�n�ͥ�n���9s{�Q�|%P�7<��*m����v����L(A�vU��"y�F�u��pq	�:�JO,��1�]+yJB��Nz��U)n`���(����u�뮈�,�x���*��
�Q}==s���d
v.Ҏ�sB�F*X�n��X�� ќ�/ي ��[3�1��9�^����r�I�v=g.�ۑ��N��-��Qu�x�֑[�G�h\)�ɽy�Oc���K�<�EE�hmǵ�l�j����6��nu��y!}����6���[3I9��)WKN��&GH�T��eӕ.�-!��s�ʳ����L�XJ��K�Q|�Ub`�ɹ��#4�X�0Ӥ�Fk��(	xof�_`�%�p2�ː�C�Е��ٻ��9Rଵ�X⒐�tۛ���i�M��F͑U�s�$-�n1�nm�:ݺ��2�l��`cE��T�]gv0$�mЊ�0q����d��j�R��jo�:]�j������Cu��	䉹~&�{�3.��Q
�y:��/�X���-�Zz|��n����YǮ��:����U��	R��ͪ�Z�M�r�c��/ԔV �v��c,�ٞ�+@B7�7�Ux�%�ǗA�	��j��0�?{=�����U�/�'�l��P���k���1��d@#HY���q��¿F�~�⟣�ܤǠT:�&7�m*ɻ��\rUZ�_n\F}O:N���d2���۝�s��*�{xt����^�`L�2V�N�x@��kEØ=��C�����]��=B��rKy0P5���;�����ϱÛ�J�F�M�C��r�z�<x@����I�8_����{=컰�ַ>nV�9
Cg��D|��2^�b�@�<k_@&귯-�驵�H��Z��qi���h�ugr<n�kz�����GY�dۣ�.�il������)ʛ��Ѳ	���vv�v��`፱�h�v�5�k!TI#�&�ܯ7�3����#�n�]��#���6h�]{�M��2���l ��x�n&��G��k�}���l�&z��|I'���m�ǵ�D&��zO�A)I�����76�Z��O�w�\$�s�YqW�}���75�x�e븑'ȥ�?���MΎxV[)��;��{�~�bvi�-��l����ƙDU������5��L)��C���Lܶs��O���z���rV�gW�K�?DJ]t:�UPX��!�l�L���(��x��B�ٝjUu���bt`薪��J�)���� E�V���.��R~�I$ +y��Wͻ6gd�$�V*p ��?�i�{�c5Լ&�B��tݠ �����k*uY��|P$�7�;�wz/�ՠ"%��\8��֫"�n��4�xc�L2�d��A�MϷ��Mkg���2"STmh	���͝�K���z�<>���]n��־ܤ��C�a��e|�|C��ʭ�h��m�o3ge�9���
&���x`]�F��f}lBS�%P�����r`p$����M��5�Q8���L�/c���frM��$;��:�/G�}M��O7*����d�bj�K�����ju��Ug+#$η=������i����8k9�j�����]��H��;!�򔲁�>���p{���k�@�����%�)�ψ@���{�g���\�շ����,�o<N�&*�u��.}9�S,O�sf����8�aUr���Ν�"]����ggF�������7�gx�EK{���A��z�����+@ZTX킒K�ґ~J�����հ3��΁�~?a��2�S���'w�a�� �l���ߦ��-T�Y��<7oMr�Gh)gn�>c���~Ik]5Z)fZ������qif�i�7��cz �d�X<�8K��L��@��,�*�=6/i�qi�����7��|��ƾ'#")^��F�R���G������uleV�GtT�M�r�v�����1��;&:�u��B.��F�h�y�)�z�z�?A���E(Q{ŉ�8`�KP�v���&�vZdv���.��_�Z�v�՘�F7P�7�g	��m=��9oZ��Noݐ�޻4�A �ۓ���	�$���������V7�WFI
 Tgӝ���٭:���Z�
��j�n|���hҁԚIў�|���i�)oc��yC�9ϲ(y(�\��Ѻ�o߈J&a�H�`v�^CJ��<~���R�!����0s`�������8<3��Ҫ>��G��OiV�=R��9(yv��;h(�*cg��P� Bצ��{q n��Ź0���4ʂ�H��1G�̉�`;��6NrdA5#;���Y��w�2�lͷ��y�n�F�JSD��p,{�l)k�w����Ȳ��>,�<-�=��A�/{~}R�U����w^It7s�T~��G�5���E)UiaSM������������8*!ɬ��E] ��@��x�z�<\�7Y��{U�6w݊}��C/�m,����fT�����ao={k7�;�Em�k�6�U��'�:	��6� [B�7�.��Ϻ�i�n����C��n�b@�y�w���o{3�|�ƕUb�7�o����-���̶�s�j�u�[q����y�~j���wL3�~A�����ۯ!�Ug��āu��C���	Z ���0l!I�l�<��[>ۏd��dֈ??���Y-��y��c����c�߅�,�OP����w�{Y���O_���q55%��~�0���<�6�1�	GU#���c�'SC��&$S�$1�9&d{ų�upRp�E+(H�R�P�����WN�iZ��ҽp�ĢJ�H=�/'�;:�^Ϟ�n�i�f��&#6b��of}'u%�%c����P��C���D-uP��I����p@��K}��͞������ ��v>^{<E1��r��b*��#x-e�z���ɉ���X��1��Jcc8��5�$;_��s���8}��m,���n�W�r߽�/����sQ�o��_y��7��}���!�vtwc��j�pY��ڭ'�[;n��Ӛ^P��.�csQ��ʔV��;NӇ6n�E�N(��C��g).�:!��YEtMV�g��l�l��Ho7ۙ#6W��T�3�A�{�^Gg�Q����C���'�4�|�4�ԩw���2�ʜQ�lV�i��z���1�˺^�4�&���>�����p�<�����uO���m��Ns��{�VG�%fg�t;s|���珕��Դ�M��ݬ�y��k�_k>���
��2K�������oiK�����`h�z��j�r5�'g,�*�N��7+[s��Ǉ-��cl!��nlrg����ՔV�hָMsx7f��X�wY���q����c�N �!f.^�cñf���8溄���4���70q(یv�跥�փ.��L���+c�v�˭��ϩ��{:��ꮫD�#�d�Rm�w.���ŉ�ީ��� ��˙�b�1Q��z�<u��6j��큻nvs�o'Y{�����%��m��:���ZR۟ң�{Hc��f#D�����u�d�qk�+��u�(7;��湌X��p�,볲�;/=
a��������؛C�<���f���m���s�j�}�����v{r�1ۋ��b�k9�#tn��!B���1����ԕFw�ny���6^Q�����*6��O;�Ɠ����"jp.fU�OEcN�C}gX�0��
ր�\M݉�V�q�YQ�X+I$ e����Ӱ��鸟'��C!6�>Iԉ�wםY�z�&��-��`�����L��)ݧ��;X�2`%�"�
y.JO` �.�5�$�˥���B���B�Y
�H� �l�h!H>��x+��f�tq"iA5�: �L�r�-�P��I�ɷF|�T�۾�}�I��S�V�R�k�-%�a���唵��w0�(��Ԡ�g��Hv��Ëw$N�n�F�c�U-�v�*ʜ�2��D\/nඣ��b<$칵�1��ӊ5#)B���Z�r=�6-��ѷͰ�pر�5�G[q����*��cl��ɍ���'g��i�9��.5�ܳvC�K��fM2QYH����b���\�n�iWԌ��D�b�5�6�ri:T�Z�?s��!�	�&��Tߧ��Z��a?5&��03M��f9��j���mvMnNЙH_<"	;�/Iq���&��|���"3rq+�/nM����'4|���&�4��{�C��� %|�*��)Z�)"�v��m�2"I�(��n����.|Y�z��D&������+���
��(GY�*w��B�A��{��ϐ���l�,&KfXp����#�.,ƶu�������Nn�=�!��Ԅ���O^��7�CGR�% ��~�S��?V�g���)I�F�Z�!6���w�{JsӜ�R�إRɂ"Q�uXX�	]�xm+	�̨�Y�:��6��L�����O�
�F�!�$���4��,�6_m�^�xB�k�i��,E�E�z=��� �:ۖ��3w,YH=ݷ�ndD-1N!{3�8�6�潖��vT���=�=n�g,c8�U�y����qp��/?�b�z���䞞u/��o�y�6��� ��X��Tti��Nv�t����ժ�<���XQއ��3�����UQ&��σe��b�A&o5��1�A9o 	��5�;����:��.y��ϼ�D�P�iLw�<��P߷�d�Ȁ�|wn�΃N�d��N�'[ʡ�Osob�%hP�Y�Z���X6�F�Sw>�����NUj��{���5ɜ�߃^�i�&`Ԉ���E$x�uWP��QeZ�P���i��^.�C��gx��L`ogs�)X��?����{���Qk�'�þ���9Z�ּ��.x38u�M>P��p鼓#��4o$=E& �r�_�Gě��H���L�C����K��ܾ����T��W[c��n����>By�p���2��9�6�5gg�b6�;ss�nt6�Dn3d�8�]�I��S vׂ�x�����뷅��/<=�t=����S�\vz۟����1�Գk�\�ڃ3-�*��<��!��Jf��σz�[6���"�vc���%�6d���u����:Q��'M���!H�s�T��'����e�hP-�ռxCO�S��Έ�DUo?3���/�A7ζs���M�j�ą�i�2M�3��7�|C��uG<�y�O��qT��ŕ[B�!�6nf�y��AQ5��~�ݾ���-w$��f��Zt�M�n�>����U~n���8,qi_��(�?}�YP�ueQ���۷V��;kD������2��,�.�ӛ���GVj�ì� 7q�m�Ǆ���@�̛��U����q�}z���P�V�W���إ�}<ĚxN��߆�׃��>\3"���jt �G�4�"XZBE�"��Xi%����M'J�y���l�p��<܄({AD�>�_R,�ϑ;�oZ��9Ċ���Ae�U�sm�/�P���dHM�u�a,��~�=T��Ι�����e���/C�~�A�Qz9N�)��4��hj p�l���Ik�4�� ��v������"���g'��6z�U��P�MOI�K��\�$=�5d.=�f����������81�.�f��U���v�3���ّG��T���xB��ӴR
o^�ȻC׻'5'i���6Ӝ3�ar���L��ß�3���w��q?�inKy͌���:0پCSs���������1�c����ۈ�^ɾ�ZbUFY���h|�J;��
$�0����oQB��N��.i=�$����V&�n�҉�*�"��m�s�="�t��S~���D��>�k����z>���t���q�^ I��{�W����d9ؽ])=	��rw�᦭�!��S#�!�I���JJz��O=c�kgZ&��/g�.�����}P�=[=V��y��](�ڍ��X�:}�l����$	ۙ�k5�GOZ�;��&-/����6������lnzݴڋ��l�U��vM��ex;H[nǖ�<v�Fm�l�׮�׆0�mNr�([�_�5E%3j}x��nL�QQ�m4�IGm�$V�im�2�\��Ks��Y���V� ����".\����SiEo��>��V�ٜ^M��FdP/�Q$�ԝ~!�,�,���
]���{�^IĆP�����o��kY�=\I9��C^��7�����:�Y,f!dp�A�Ew���҂�3��ֻ8�gR����um���RK$y|��^�W�.*�� a�w�H�1��%��� Q
2�S�T(?Y�װ�k����:p����وNScOS�/#s--��I)�#�n������+6:�J=k�W�<���ȡ��֧}�����5�xv�i-D�s=�;����ˡ�pz�wA�h���m��
�t#�p�uE ;5��ö;�!�׽Uy�z�,������GhkO��1S��>!��[TßCU���\�Af�85+05HĈ�G�)Jܙ8ݙ��ܴ��p��z��8!�B.v�<f*��u��ێ�{��"����ӉU��'������G��r�R+2���u�y�28�l4�����{��E�q�U�~(z\�k=g6G%Ӻ�U;y� ��B�U�A-l���Ui��L͆V9~��Xĵ�f[';�l�yWdE�I�]ۙH'���V�R�q�μ�ӗ��wt�Y���{���T�;�{����|�5��G,ĭW�?�����	��n�ej���p���=ѝĚ\��|j��6v�a��w,�t�3)�mG�ė�<��O��w�_ c��]{Lz�>�8�����U	ډJ�n��}��\�X8�1ϰ�hu�Ė���=n$�=N���.RZ�bW�r/���<6t�s_\�Y��.�wG)1�t�ͱ}����{�U�[���b�[�p5�ھ.���fV=YS��AD�˳��}�sw:�涝mq�r �N��61p�a��լ�W��7}Ns�}T��{�i\=��e
ґe5ynU�-ٜzCU�ytvA�o�L�����8�gp�PF����p�8\�Zޭ���Wxڗs��&�GD��`9W�	v.��P���5�6X�A��-
}���ݼ��:�\����������\�[E=� ��x����y�EE؈]��ئ���s)�u����"lN�yY����~��n�Vl���$>�l��i�U�\��ui��E���`�J�̘��=���6�C��Kl 1���MX9k��"�����vml�ST>�Zyi�֎z�Z>��cڤ���3"��R"��{�ȹw{��5��U��>܅��v��ޤ�̊iTTB��<w�}���%Yl��rev�����sgy��X�M����
����Y�&|̰��\:�nuZ��A_E����DAUG��>G�Z~��ހ�N}Z@D6��p�Z��2\�݅�-Ԑ�IL�L!>��g��n���M�y��
�꽍���?��ï��+~)A�{[3O>P���oeսg�,��7��ĚLH+�>jL�)�E:�Ho}�q�����ߖ\�����Vu}�\�I���g�'DЕ^�AZ�����*v�D���X@�͖� �I��Tdn��� ��q��8�kD�;ZJd�w5�Z�.{O]nq��n�������̓�FGs�6����uk-����t��s]�~��2�C��;�r�ݦ$&���o,��I&�h+�Z�\&�-B�W/{��x��t6�[�G�yp���W�R�=��:��̋�E*-��ތ��*}��笖��{$ޤ�^�]��Ow5��CU��SU��c�A�b$���{ӽ�P5�t|c�+�����g����5,r�Z�l��Q�(5Z�u����������Z ��Fo�<�f�g^����y?���Ң�,�Pj[�`,̕3�s�����w��_�<�A �gL|T+��}w�3��?�L��jh�����iOxC�P�4y:[u�,?�?j�3��ᭀ:۴O�pH�'<�>�
D���ɯN]l���h���hr$!RA���M�2��m�g*�PFh�#)�S��|�[��\5�	�'������n�B����	�g�s^��[�^�[�%,39)r�V ^_u��:u��U��@D��Ə�iu�&�i��ڲ2(v�` �4�+av�����D]�f掹DW�c0m�g;G�n�Sq����ߺv�hȢl����a�<ǟ��u�k�^j�
�	�Z�u�ⲏl�����u9�t.Ó���t��M;Y�v�����!�F�!��ڜ�U���<O�@�m�m@�3�R^)��>g��B�����T�X�V�y��]��!D6
S�.21l�Q���(_QO�k��9�D�-{��>�͒^P��i9�g���p_�v0�N�~�L����xY�lηc+�{�
��UY\dq�V����|,�j&MD	U��W�3+���K����h��>��iP��L�������{H^�

'S� 0�m�S��!zꢘ�zM�C2.�T�e#C��~DUytc�'��K#��e�{����MP��\hQ�����JX�\VDZ��x��j��R�qV䗵ن�/ְS�\ݶ�^�e�<F�h8�vz�G��x�wg�ONY��Z��ݮ{VN��GE1�)��G���7���"*'�n�}�.!e����(�6�ub�ϲz��uųͷ�1�{!��D��E��ʻ@i����1[{��)eP>��Y&߾�h�����Y	�7H,��� �6w[�W�D7U������}7������!�ij������\��k�KY̌܇�8^��)��	-���»�%������+O�M^[�"<6�����y��3��pK}�U�ĺ�����_
k� J�\jf�?<�S��M!gi�;��^�����L9���tб�C�q������JeP_����p��i��U�쓻�����bM�#��5&�
����v�3{d�.��(.�T����ak��npv�1���U0H�3ˆ�B�R�ϵ\��� i���(
�Z�/�ӄ:[5����H�	NrYEOt}��Đ�
�y�����}/���&��g�	�QdU��0�)eH�nP�u3�/�j����i��*�T�8���[+����C�>?UJ9W���P��4���9�-��+���hxW�{���c����Z���0�2�oi,�F�-.}���/{�,cMV�PO�IH������^���r�"�b��}�����oǅ/2I��=uP�j�^�Q�ް|�H|k�����e�Ə���G
 �`� ��p�eFx+;M@ީ�k"��-�y-Cy�07��em�2-��xK���;������	F�J��uW�;V�5����	�|�r�����u�T�ם�ft��oV-窣$ݹ��{HZE%���8Xk���N�m$-[��ˆ�Ȃ���_b�)}�^ٲ�x���;�D)7�uY��������q�Uky=�Z�֪5��J�()��X�)o��EZ[Ț�{��>R���UV*��aj�Xv,eND�SMVR���c{��YZ��nuv���xt�Z�ȭ���-���0}�xl�wA�I���ξ�f�nR�5L.dL��{�]��ppR�ׄ�N�x �<���u1�������7�Ծ޷�̘�G��.���vU���L�iv1�5�al�e�o�%�ǰ�+z<�p���^���߆V��h�gE
���憔���c���(��[���U�}A+Ϻ\Ml�k�������m팭���r�j���$�F�y���+���:�ގ�0�3j���[O�{�����ؽJ��B��Bk,��J4�0��f�9�S�ce���Z�g��uPb��n��k\�]\�M�ͨU����\�\b�=$9�&Ev�wg�f�3�������<��b��n9�CqĳƄ��B�]��y�۸���w�S��ۆݛ�v��pNի7;�ط"翕~֏n��)[�"�:|��{�:��㍮ޘy���6=6�b�`�ζ�=�+��ut����r��=3^Tn��糱�<��<�������=^��Y疛���u�;u�O7e�.��bo=r�b��|h��8t�Q�u�D���T��%���p(���<󫮓u�V|�n�q�t�a�.x��ool[h�͐�n�\������ې��9��e%o:��S#�t�����|��Ss�m�ێ����Z��\���`��\�9���p��q�w�rn>���ٞ8��mŐ��2�C���C�.'!l���󬴑���u��MU��Y!��;�vu��Zۮ˙�)w&�#��0t��s^�:����+E��Eu�60��hoP]{a0u�Z]	z�32�*2sǅ`��
ژ��L�{4F���\�a�IF��ym�K��pe��>z/�kuw�37G�}p�K�����h	h2l�;-�׆�*�p�],洙ޙn��8bUK���n+Z��nn1��h�qYSn�a:����r�Y��_c��	��f��:� ���]e�1
<�����1<ї�&a�Z��6��'<׉Y=]s��W�`:�����6M$\�c�z6����V��G� ���ݤ��tĜ��w�y����::�T��.�npNz�U׵�`�'�p�l�$�nv'��K��bؼI�̭���ĉ6��(����)Sbw$�Ś��H�߷�=� ��������|�"23B��z~$|;��������� �qG!�a������#9�6�h|'T��5�E�
s�(A�2��+�6P΋;�nY����R)_[�Y��Gl1���ͼ5���|��׸��P�d���j��ȼ���	/5��g�J7ک�e�uz>�abf�L�k����^�e�c�]��_���ѽ����yE\C3��;�3��ẃ��� Y��a�����*�O]z�pX�����^�`���"}t��,)�-�U|m�y�W����]�� Ԁ���]�i�]�U�W6mn
�ױ�؞N�>�mz�fOb߁U�g�uH?"}��Pbb"~�Wu?��`+r �tb���$i����q_|�*�uF�!;Oݧ�հ���!����D{�;ܞ��I3� G�9M�y^�~����`I�n����ylw�J��e�N	�)�	� �lR�+�	�ҍ����s��0%{7��qV�w�>�^��M�~��߰B��k>n��m�y���)�o��ϟ����޶Q��2;��o�r�g'�,�ه"����.j�M�l�KY��}8�a\�	M*=Ąʜ�D%��|��[���rxlC�E%թn)iGe��JG}Ń:jkJ�9{rgq��E�*��?v ���׌(s{�� V/��&sP �^��]�R�b�
?���Rw�PT���*yWо����q+�c���
��x�:/zi��#�������O�b��!ʫyv��G?�7\���Z��9�M�鵢؛WI�U�� �1��f����P[�`O'K�6,��t���e-��.ښα� �����TW<࿑H2Sd����[�!��W*��O�Oa�4Gb�tg�Z9���1�f�n;mMZ��l/Sw��6�s��|�ת[�������Y�%7�RK>�Շw���{���˛���a(f޼�;�Ʈ�sZ<�W[���e.�[�Lq�5�~HU|xa���.w$�Qnz�Ά�;���޶�O�{�_sN3~U({�0�}��q�Hk�����34��gc.W��ܿ]�?Qo,T��o�xK�f���DҐ��ݑ{�E@�"!۹0~�D{�D}if��~�$��2>��6���H��U�w��}�X^��Np�{�҅ @��Ꜳ�0z�?�U����׸%kK�Ʉ�K`��;b�2EW��vo��ݨ]/N�������B͂�'���?� �2S��T!����&��Q>�P�$�7��H]� �L���M֑Z�;�cuq����}s��3k��,ǲc��X��"��c �c�	��̄�#M��}��6�����w+��X�Ƴ�|N����g����
U�-��s�7��4�7�t���W���>�Z���pw��D�hAr=�R�Ҁc��y|����8L+���赴�m���z�x(��������J�ׂu��+�M�Q�w�Iw��M���W��e�~��<Au4<��鬰�vY�
�;y���vD:ڈ���~b��<���DOՋ��W�Cә�o?{dO�"�;��� �eLu�u���Y��2��<���k�+�ӓ5���Ǯc�B��3��a��P�pB����p>�����j��v�K1뚗�U!W|��myeK���*�KԆj�5�"J�1��-;qh]9�k�k����ŝ�~L��h��x՟��<<xƱ�cq�	%�n��f��uv:^�cu�����.�=M�^�=1������Gd�ks�PԀ�m�0�Y������(jq֞q�ސ;�o{W��^s�7�6x�8�k��B����L��DIP��)��� ��ezN{ʜ�lj�n*��W�|;c�[��(Y�o%0@�7���y��Ps��>Ք��0|p�J2��K���^[hA]�>�]�o�A��8�-x��)T,Et
XBw�&�oXT���)I__����q�,Ϸ�9I�H��U`Y�#�"\��4h�@�"-S��mW�hjC�;{��S3���"n��[Q��y&e�a�X
����TY$���\����3���0ßu��ijE@�F�����|V'�����}۩�������1�����*��o�x�z�=�F� qJEZl�-�[���`k��֩�X�m��77g�S\�Y�7�K5��R��E��{h�k���jkʥ0D\h�v�����Kf�ʍ���a���]W4V�DX���N�L��r��ܭ�Dl�|y��-T�NJҮT+�V�ùh�tW�;���n���:e�Ƽ�'��I�C5��X��Į�^�*㘁t�@rr�W�{�r(qл"6\��7)K�I��/a&"K��w9T��gn��ۏ ��;��:o2g7;;R�w� ��=�Ɵ��L������A��=�Q��w��iמ�M���y{4|m���Y�i�N��78͌�s��6�]��X�n�)%��sZX'�]^N8�/�=g�3�-(ӄ9�g%��o���1�b��q�������"opOV(��:���1������+����S��KHA;s���\_6p���yM)7+�m�2"7���B;'�r�����3j`u�8÷�;ʂ�<�MJs(b�g��f�!�fX�X�M��ga����B�[*��[o�o0h��\�Y��0�g62�gHѣZݚY�N'�0��X3.��X&X{��,GKx��Ӽ���r�gl7ofp$�.�t���{ܲRg%��pS0�*�[������4�E��ɛ\�u���c��S~;s��ڹg�)����Gw3P޸�������ռ]	(����
W��GRSb� ���Yd�䆧rw�K.��av�{ѹ����O��H������F�9�*�w�uqgav
�������^�ʹ������Ɛn� p�b�Qu�Z1
'�@{��ШD��_kJG���Qak�>��������-UBTP�+�HGQ*�ZDI,�ugs>�3=�Ԡ����=g�]��szS{�,��� gڅ^���ym��m�$^���)Ly�NM�M��T�Z���� �=��*��\R�ֺP�v�fT��JVyl&��r�c|hlw8��[S}�ʣ��m�:�=׽�u@jy���+�rU$���2g4%�ގ�֚�}IJ��Iռ�P�oXa�GJ[NLӗ�
B9����p�Y���Eo����7� �S5lz��uG�cĕ5��(�f<�T�yf�y��Y�UM�47�Pj��婶h��+_lO޴��ƀhl�K.�7��c�&땂��ϵ	�ٻ���n���v��N'J�ڮq�^x=�啋���e:�V�M�u�ݘ�\��R�8��5n{4���9�wR�NڵF(��� �\�A8��@����K�۬M/�w����b2��Yܼ��w��r�snrֽ�	Լ}��WΖ3��K5�so�Us
a?e-ID58@�+�=������Bw�0Y����Ny�o\�`��E؝�"�"�b�H�!� ��q�Dm��n����gzqr���s�7M'mp^�v��n]K��,z���IaSu�=�0�C7��Vh�:�yø2wׂIƦ<���]IiQ����'HU���z�a�*s�M�Vξ+�@΀G��cu9U�?}��8�z�L�~]���L�/�M���E�D7�#4&	�V�ծJ�4&U��~�WG��W�t�m�w��w/[��HU{k1�o�����p(����f�,e����=�2E�lX�b2��x�"��>�,��P2J�-�F��ɢ�8m��Oш�&$�U6���"��;��s�t׹��π ���yH��a�&��-C[���9K}{ƾ�漱���o���u��n��`-,HeeJ��ߦM�� m.�b�b>s~\��r�'��f��B���p�a_z�JT|�gھƢ׏��3њ)��g?�pF�>� �217�8vF�;.��c-c�9��񂟉YB�l�)�ll��J�n3S���>��F�Ilg�{�3
n/��b��d��)c����
UeQ0n�kY�f9s���^�n���C�if}X]-y�Oǎ+)��w�e]���վ׊N
��{��c��o^I\ǳ���ľW�v����\ƽE.�-�f���� W����7�����m�o�4�f�{����'��X��Gx��z�T�4V��u�Mұ�=lv2k�vxzs��ٻv�;���.u��tI���s��ݻ��g[�x�][�vp��氽D�u\���"��f�v�yb�	ɍg#ksi�k�-o�7�Mu� $�J�������~I�/&k.r�{7����9�r!1k�>x�K��DЂ#���n~@J"~jr�s�~~(�kl�F�ڣbX`�nc6�W�������4��
��4���8���0B 2�n�%��F��]�%r<�&}���Ϥ�`�3W���:�Z���6'���S�_n[�B7cD�c5� �A�H/��B�j�ef�QI
uB�����w.�^g����)� �5�=0�K�a?��P��i~�����;�����e���_m)>)y� ��o�QK��F��]ƃ�[jKj�.�"�ڶ(p]d@uM*�}j�{�D�מ6rz㹬0��\�y���ꄯ��X	��(��wk����#ǖ��#���a�ٳ��H�"Q�w�K~K���бm�j�+�oX9ć����G8b��B+M��4.��3�>����^ {�z�
l�J�Ȍ�!��gL��ۛK��/��U"�*�Ta�0�EW� D��;�]���0>�U�[�10Gf���KֶUA�`yt<Q����` ғ̯	�u��dy'T����ŽO/�ZkpV8`�$�/����Ã�U�.��r�=\�w�>[2/��/%�n��fO��X"�	�?+biwo6������y; �uPu%Q6�h{�H�y�r��yE'��:x���R9W�H~��	��1�ި<�}��I��R��:�|k�q
'Aؾj9P�uU{c�
�Aw��+WH���y~��U~J�ШJ�޿Z�4�n-��UU���4�ͳr���&�f�~��-��Y��pV��*�[�(��؅�����]�Oq�.77L3m,�3K�,f��m�l͔f2�3��EVcu��4bM��n�s��t��Nv�;7lv�lV��[p�۔�3�퍶�q80�3m�Y��˙����<m�aˉ�m�n�����C�Y����g:7;�q�����������zs���m�jͶ��XUSx����8�WK���Ϟ|;~��?��q�^,�߾o_��z?��=���]���.�w�.��o�����_������O,w�<�-�o�������n>/^�s��WMۺ�fٿ~=�ׯ|�׈�o�~��Mɾ�ٽ�2�lm��Ŧ�m�ܛ�ɾI�ݿ�Ӻ����L}X�v�7!o�ǣv����߽���t���Y����X��?;m��}���{?N��쾝�������<-l�n[���};�g����[AѦX�|Nw.�~�Tpp����[���vn��n�\�ۺnݮ���|������7N3��q���;5�>�忾�x-�:ݻ�㌲��YE�2�E��&�Yl�"Ȉ�ȋ,��k&�"i��k$DZ�DYdF��Me�Qk,��D��ֶ���&�"�Md"�,��Z&��4[Y4Bki�kY4Z,Yh�Z-�B",E�[,�-��Ybɬ�Me�&�BɢȄ[D��$Me�Zɑ4Ydֈ�[DY"�k,�Y-"�-d��h��ȶ�YdE���k$Ye�D"�md�,���ɢZɢ,�D�K")��&�"�h�"�",�ZȲZȵ�5-dDYe��d�k$Z,��YdX��,�"�B,�"�-�,�DD��Ȉ�,�,�,�ZȋE���,��i�k""�Z��DE��YY��h�e�Ye��,�Z�DD�H��ȵ�Z-YdMe�Ȭ�$Z,�Y"�,�4�e�D"��"Ŗ�h��+-E��"ȲȚ�-h��Zj-���Z�Z%�(��-4���D��DYe�Ȳ&�k$Z%�,�k-Ym�h���D����K-�ZDY"YdDZ���DZ�Ed�L�H���"!e�&E���E�E���Z�,�5��$Z%�DYdB(�,�,�j%��֊��DEdE��M�D[,�,�Z��"�H�Q"�Z�%�EdE��Md+E��k�D�DM"h��k!�֑me�X��eb��Yȉ�L�[D�e�YD�ȑ,�"D��H�YE��"MEe[K$Z�h�Z+-,��YE��VQm4��e�YZ�5�-�%�idD�Y"�$M5H����(����VimQ,��"���H�K++5j+%�,��,�j%�V�d�E���"��$VkD�e�"Y"�K"��Z�-VQX�Y��mb�iZ�X�,QYEf�%�f��Yh�M"�d-dY��-��X��%�d�b�&K5�Eeb�)��ڲ�+%*��RE5+U+U*JV��իZ��MZ�j�V���VVKV�J���e%VU)*KZ�j�Z�~瓚��j����U�UjQF��[V��Jի2�5P�MEPE�l��ĵ6�Jj���Zn-�j�e�MIf��$K(��mEj��+$Z���:�ny�%���L�H��$S�����KQ4H��-d��E���mYX�&��-�Z�"��5�E4��-�Yh��e�5��dVY)��b��e���(�e��D-��X����6�,�h�-iYh���E�-eh�[Z�Y0�YdYe�ZYh�-��EdD"ɤQb"#k-��k",�e�Ed��"ȵ����D�,&���ڋYK,�h����-5�,���%���ȄE��"�"-e�H�ȈE��D�h�5��D�5��kuոn�(��e�!"�YE�k&���B-������h�k"ȶ��,��"��D�B-���D,��Y4[E�H��ɦE�h�X�b�h��h�"ɢk[,�-��F�,����!�h�Y��kE��D�"�"��h���"��5�Zh��dB�h�MdBȋ�����B",Y2-�l�[D�["h��D-i�,��&��-�X���L�,�B!dh�ɢ�k,�����i��Bɑe�Zȅ�E��"�,���DBֲdX�e��4[Mb&�h�Ŗ�k&�dMd���[Ym,�-�-�f��M�D�L����dF��D�B��me�j&�Y�-���l��M�h���"в�,E��!e�F���[D"h���,E�&�dY���L�l�e����m"e����d&��M",�B,Y4M4"dX�ȶY5��5�D�X��ŵ�Yd�e�d�2#Y4X��Ym5���dE��,�-��ɑMd�Ah��h�e�X�Dȱ4�dMe�&Y2,Dk-�h��h����-���-b&�h�e5�L�"Z,�"&�h�,DE�DDK!,�Ye�L�YmZɭ�i�DY2�D�E�E�"�[Y2�"E�BkE�M�Z"-�����m5�E��&�k-dȚ�Y2-�ŖD�Z&E��Z,�ȵ����-���h��e��L��,�����"""�M��h�e�",�֋k-Y4Z!d�E��YdMd�К�����r��lpw6��n峅�o��ܭ��w�o�x7F��lm�Ÿ٭��-�۴uo��7W_n�Xt7;q�~�Ѽ;���&���<v���^�Vv�����F��F8xC���ߡ^��o�}���{��nc��nN��s�s�Y����]���o~�c�vo-�C~�ݎ����zz��ݳ}���7�۽����7Ѻ�t߯&���Ҿl}�������'ͷٽM�m��o�����.q������ǥw�wnﻻ~�{�[�{��oS��w�޾�W;m�l�[��m��~������O����o��>�a�[�=-�w�Gsv��;��Ѹ1�����u=aя$�n[��8ߩ幝��1��fCNɺow��3v:�5���������MÍ�ڶ��O�v�;v�i�v����q�q��t�:n��]�8�;�4��?S���7�q��w����f�A~������m��o���1՟���{�������9���q�>[忱�������;۽�Ϸf���~�ˆ�C{<��>g��o���x�Λۿ3t}տ+z��x�v7�i��٭���y�o�-��߭���f�o��ݛ�n�}�;���V鼶�ǣ�oͻ���۩mc�q��O�ͽ�˦����5��m�kz���,v���?��oI$�q��c>�徽��۸u��Jy������cz��O�|<�����٦~�F�7��m�φ��h�9�w�SX��ǹ��F�#ug��y�k[�Cww{=z|w���O��r��kv>m�q�{��A�M7�����>v�6��]��o[ll�o�r}�ݼ��83����h����a������޽�Mٞ����~]����3{�K�n�}����ǳ��q����7��m��ն��]��BC��8