BZh91AY&SY.�� �_�Py���߰����`����"  ��m�G M�Je2'�FMOL���hhd F���%FOP   d   � �`�2��Jz�&�D� ��`�	�0&E)�M<����� @ �"A4&��I�z�<Ҙ�"h��OQ��%
�V�����Q��(����=���-Hb�" %*W�G��,�Q��6I�����4�ʀ4�u��@x�e5W��"�,��	DI ƽ���1N��BJKy�*��/Ii��Pc��n�r�&
!�Et,���3���b���"N!��h=��j)�Ǫ"7r>����͆!R%����x�þ;��¢͵{�Y�g-�Q�na�r����)�܆�"9,�`�Xlek4! �Vq}B�4-#��߆/��zI �&6?:�|b���8����&�s���K�K�A��ܯ�j̥VގH9d� ń��th��zY�3���ԺǏ�5���p���SK�y�z��'�̦F�i^d8�8��Bd[
 M����l:ڞV�a���r��<�(�E�0y�<�Am(m�^B�G�2@���ll�@�#�F��;K	��X�l)
���SO$f*\����&�.:��Z��4�3u	f��;Zvl'پ0kx��}�iݶ�Y��Rw\ڡ����ùQ@��[;w̋���H`؈S,���lY���6��u'h^F�!��On��0�lU^���䖊ETÇa�T`�|�(��zˑ�C������VH���ؠ^&w��
8�$��L��>%��
C�<�N�bE��AP�Y ���M�#���Y�"�wE8�c҅��1�g}�]rEc���(����EWfj-��a�ƙv��N�e��k-gM���iq�"�V�<Sb��K����{x*��ͷ�m�+W��i�.���B �PAZ��^	,��Pa�#j�Е@����#��ؗD;5�9�r(�&I,�v��y�eTR�I�!!B�cA�R��^�4�L)�
������` cTa��H��K���u���\��W���~��h�T�8�3�8���R֛U[�Y�F7Ⱥg#��$udbIm�|��\d ��z˕X�`�����$���}�h��j�w
�<��P��a�\�Jw��(��3<5>�G������W�~#lTD\(Z2#�F"�C�a��2"�%%��X�$��a��4B#��z�ۃ�e�u�>��td�]V�*՚m�2��@&��PŠ��N���(D��@����v��]i$$V(�W���0�.�ԼfoN�ICZ���&PSg���v{�����w� �%+���F(s��9Rx�T�9��Ē��&�������͠`����P�7`�m��D;׊RH
f���=[���R9��_}מ���h��^� �I$�̽]/��:� \ �`�]�����1�dL� �� �F2�D���� &Io��I
tCN��5$����}P���WD�B�A9�pRL,���*i�˲��dN�@WՐ��쁩%R�,=-flц�Ɍ�Pp�;�΁�"▜6S_�	p#F7mʺ�Š"�[�.���7����|��0=j b��
��D�i�A dA$�<)G&P4S:N{2KU�J���eJ�RU	���v;�I ,y����F���3!�cJZ�nS��>�6�<E�G��L(�����v��6$���G2GhH�b_���X�U$�Z�"�8q�W�Z���ײ����'�gi�2�(��o�]��B@�`J�